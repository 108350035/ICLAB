module CHIP(
  // input signals

  clk,
  rst_n,
  in_valid,
  in_valid2,
  matrix,
  matrix_size,
  i_mat_idx,
  w_mat_idx,

  // output signals

  out_valid,
  out_value 
);

input clk, rst_n;
input in_valid, in_valid2;
input matrix;
input [1:0] matrix_size;
input i_mat_idx, w_mat_idx;

output out_valid;
output out_value;

//input wires
wire C_clk, BUF_CLK;
wire C_rst_n;
wire C_in_valid, C_in_valid2;
wire C_matrix;
wire [1:0] C_matrix_size;
wire C_i_mat_idx;
wire C_w_mat_idx;
//output wires
wire C_out_valid;
wire C_out_value;

//core module
MMSA CORE(
	.clk(BUF_CLK),
	.rst_n(C_rst_n),
	.in_valid(C_in_valid),
	.in_valid2(C_in_valid2),
	.matrix_size(C_matrix_size),
	.i_mat_idx(C_i_mat_idx),
	.w_mat_idx(C_w_mat_idx),
	.matrix(C_matrix),
	
	.out_valid(C_out_valid),
	.out_value(C_out_value)
);

CLKBUFX20 CLKB(.A(C_clk),.Y(BUF_CLK));
PDUSDGZ I_CLK(.PAD(clk), .C(C_clk));
PDUSDGZ I_RESET(.PAD(rst_n), .C(C_rst_n));
PDUSDGZ I_VALID(.PAD(in_valid), .C(C_in_valid));
PDUSDGZ I_VALID2(.PAD(in_valid2), .C(C_in_valid2));
PDUSDGZ I_MATRIX(.PAD(matrix), .C(C_matrix));
PDUSDGZ I_I_MAT_IDX(.PAD(i_mat_idx), .C(C_i_mat_idx));
PDUSDGZ I_W_MAT_IDX(.PAD(w_mat_idx), .C(C_w_mat_idx));
PDUSDGZ I_MATRIX_SIZE_0(.PAD(matrix_size[0]), .C(C_matrix_size[0]));
PDUSDGZ I_MATRIX_SIZE_1(.PAD(matrix_size[1]), .C(C_matrix_size[1]));


PDU16SDGZ O_VALID(.OEN(1'b0), .I(C_out_valid), .PAD(out_valid), .C());
PDU16SDGZ O_VALUE(.OEN(1'b0), .I(C_out_value), .PAD(out_value), .C());



//I/O power 3.3V 8 pads  (DVDD + DGND)
PVDD2DGZ VDDP0 ();
PVSS2DGZ GNDP0 ();
PVDD2DGZ VDDP1 ();
PVSS2DGZ GNDP1 ();
PVDD2DGZ VDDP2 ();
PVSS2DGZ GNDP2 ();
PVDD2DGZ VDDP3 ();
PVSS2DGZ GNDP3 ();
PVDD2DGZ VDDP4 ();
PVSS2DGZ GNDP4 ();
PVDD2DGZ VDDP5 ();
PVSS2DGZ GNDP5 ();
PVDD2DGZ VDDP6 ();
PVSS2DGZ GNDP6 ();
PVDD2DGZ VDDP7 ();
PVSS2DGZ GNDP7 ();





//Core poweri 1.8V 8 pads  (VDD + GND)

PVDD1DGZ VDDC0 ();
PVSS1DGZ GNDC0 ();
PVDD1DGZ VDDC1 ();
PVSS1DGZ GNDC1 ();
PVDD1DGZ VDDC2 ();
PVSS1DGZ GNDC2 ();
PVDD1DGZ VDDC3 ();
PVSS1DGZ GNDC3 ();
PVDD1DGZ VDDC4 ();
PVSS1DGZ GNDC4 ();
PVDD1DGZ VDDC5 ();
PVSS1DGZ GNDC5 ();
PVDD1DGZ VDDC6 ();
PVSS1DGZ GNDC6 ();
PVDD1DGZ VDDC7 ();
PVSS1DGZ GNDC7 ();




endmodule


/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : O-2018.06-SP1
// Date      : Tue Oct  8 16:23:25 2024
/////////////////////////////////////////////////////////////


module MMSA ( clk, rst_n, in_valid, in_valid2, matrix, matrix_size, i_mat_idx, 
        w_mat_idx, out_valid, out_value );
  input [1:0] matrix_size;
  input clk, rst_n, in_valid, in_valid2, matrix, i_mat_idx, w_mat_idx;
  output out_valid, out_value;
  wire   N942, N943, N944, N945, mem_num_4_, mem_num_2, mem_num_0,
         calout_num_0_, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041,
         N1042, N1043, N1044, N1045, N1053, N1054, N1055, N1056, N1057, N1058,
         N1059, N1060, N1085, N1086, N1087, N1088, N1089, N1162, N1163, N1164,
         N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174,
         N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184,
         N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194,
         N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204,
         N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214,
         N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224,
         N1225, N1232, N1233, N1234, N1243, N1244, N1245, N1246, N1247, N1248,
         N1249, N1250, N1251, N1252, in_weight_flag, N1276, wen_in, wen_weight,
         N1286, N1287, N1288, N1289, N1291, N1292, N1293, N1294, N1302, N1303,
         N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1321, N1330,
         N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1349,
         N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363,
         N1364, N1365, N1366, N1367, N1368, N1369, N11306, N11307, N11308,
         N11309, N11310, N11311, N11312, N11313, N11314, N11315, N11316,
         N11317, N11318, N11319, N11320, N11321, N11394, N11395, N11396,
         N11397, N11398, N11399, N11400, N11401, N11402, N11403, N11404,
         N11405, N11406, N11407, N11408, N11409, N11490, N11491, N11492,
         N11493, N11494, N11495, N11496, N11497, N11498, N11499, N11500,
         N11501, N11502, N11503, N11504, N11505, N11584, N11585, N11586,
         N11587, N11588, N11589, N11590, N11591, N11592, N11593, N11594,
         N11595, N11596, N11597, N11598, N11599, N11681, N11682, N11683,
         N11684, N11685, N11686, N11687, N11688, N11689, N11690, N11691,
         N11692, N11693, N11694, N11695, N11696, N11773, N11774, N11775,
         N11776, N11777, N11778, N11779, N11780, N11781, N11782, N11783,
         N11784, N11785, N11786, N11787, N11788, N11870, N11871, N11872,
         N11873, N11874, N11875, N11876, N11877, N11878, N11879, N11880,
         N11881, N11882, N11883, N11884, N11885, N11964, N11965, N11966,
         N11967, N11968, N11969, N11970, N11971, N11972, N11973, N11974,
         N11975, N11976, N11977, N11978, N11979, N12060, N12061, N12062,
         N12063, N12064, N12065, N12066, N12067, N12068, N12069, N12070,
         N12071, N12072, N12073, N12074, N12075, N12086, N12087, N12088,
         N12089, N12090, N12091, N12092, N12093, N12094, N12095, N12096,
         N12097, N12098, N12099, N12100, N12101, N12102, N12103, N12104,
         N12105, N12106, N12107, N12108, N12109, N12110, N12111, N12112,
         N12113, N12114, N12115, N12116, N12117, N12118, N12119, N12120,
         N12121, N12122, N12123, N12124, N12125, N12206, N12207, N12208,
         N12209, N12210, N12211, N12212, N12213, N12214, N12215, N12216,
         N12217, N12218, N12219, N12220, N12221, N12222, N12223, N12224,
         N12225, N12226, N12227, N12228, N12229, N12230, N12231, N12232,
         N12233, N12234, N12235, N12236, N12237, N12238, N12239, N12240,
         N12241, N12242, N12243, N12244, N12245, N12486, N12487, N12488,
         N12489, N12490, N12491, N12492, N12493, N12494, N12495, N12496,
         N12497, N12498, N12499, N12500, N12501, N12502, N12503, N12504,
         N12505, N12506, N12507, N12508, N12509, N12510, N12511, N12512,
         N12513, N12514, N12515, N12516, N12517, N12518, N12519, N12520,
         N12521, N12522, N12523, N12524, N12525, N12566, N12567, N12568,
         N12569, N12570, N12571, N12572, N12573, N12574, N12575, N12576,
         N12577, N12578, N12579, N12580, N12581, N12582, N12583, N12584,
         N12585, N12586, N12587, N12588, N12589, N12590, N12591, N12592,
         N12593, N12594, N12595, N12596, N12597, N12598, N12599, N12600,
         N12601, N12602, N12603, N12604, N12605, N14263, N14270, N14271,
         N14272, N14273, N14321, N14331, N14358, N14359, N14360, N14361,
         N14362, N14363, N14365, N14366, N14367, N14368, N14369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n690, n726, n727, n728, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n989, n991, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, N12485, N12484,
         N12483, N12482, N12481, N12480, N12479, N12478, N12477, N12476,
         N12475, N12474, N12473, N12472, N12471, N12470, N12469, N12468,
         N12467, N12466, N12465, N12464, N12463, N12462, N12461, N12460,
         N12459, N12458, N12457, N12456, N12455, N12454, N12453, N12452,
         N12451, N12450, N12449, N12448, N12447, N12446, N12445, N12444,
         N12443, N12442, N12441, N12440, N12439, N12438, N12437, N12436,
         N12435, N12434, N12433, N12432, N12431, N12430, N12429, N12428,
         N12427, N12426, N12425, N12424, N12423, N12422, N12421, N12420,
         N12419, N12418, N12417, N12416, N12415, N12414, N12413, N12412,
         N12411, N12410, N12409, N12408, N12407, N12406, N12405, N12404,
         N12403, N12402, N12401, N12400, N12399, N12398, N12397, N12396,
         N12395, N12394, N12393, N12392, N12391, N12390, N12389, N12388,
         N12387, N12386, N12385, N12384, N12383, N12382, N12381, N12380,
         N12379, N12378, N12377, N12376, N12375, N12374, N12373, N12372,
         N12371, N12370, N12369, N12368, N12367, N12366, N12365, N12364,
         N12363, N12362, N12361, N12360, N12359, N12358, N12357, N12356,
         N12355, N12354, N12353, N12352, N12351, N12350, N12349, N12348,
         N12347, N12346, N12345, N12344, N12343, N12342, N12341, N12340,
         N12339, N12338, N12337, N12336, N12335, N12334, N12333, N12332,
         N12331, N12330, N12329, N12328, N12327, N12326, N12325, N12324,
         N12323, N12322, N12321, N12320, N12319, N12318, N12317, N12316,
         N12315, N12314, N12313, N12312, N12311, N12310, N12309, N12308,
         N12307, N12306, N12305, N12304, N12303, N12302, N12301, N12300,
         N12299, N12298, N12297, N12296, N12295, N12294, N12293, N12292,
         N12291, N12290, N12289, N12288, N12287, N12286, N12285, N12284,
         N12283, N12282, N12281, N12280, N12279, N12278, N12277, N12276,
         N12275, N12274, N12273, N12272, N12271, N12270, N12269, N12268,
         N12267, N12266, N12265, N12264, N12263, N12262, N12261, N12260,
         N12259, N12258, N12257, N12256, N12255, N12254, N12253, N12252,
         N12251, N12250, N12249, N12248, N12247, N12246, N12205, N12204,
         N12203, N12202, N12201, N12200, N12199, N12198, N12197, N12196,
         N12195, N12194, N12193, N12192, N12191, N12190, N12189, N12188,
         N12187, N12186, N12185, N12184, N12183, N12182, N12181, N12180,
         N12179, N12178, N12177, N12176, N12175, N12174, N12173, N12172,
         N12171, N12170, N12169, N12168, N12167, N12166, N12165, N12164,
         N12163, N12162, N12161, N12160, N12159, N12158, N12157, N12156,
         N12155, N12154, N12153, N12152, N12151, N12150, N12149, N12148,
         N12147, N12146, N12145, N12144, N12143, N12142, N12141, N12140,
         N12139, N12138, N12137, N12136, N12135, N12134, N12133, N12132,
         N12131, N12130, N12129, N12128, N12127, N12126, r1350_GE_LT_GT_LE,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128;
  wire   [3:0] cs;
  wire   [2:0] ns;
  wire   [7:0] calin_cnt;
  wire   [3:0] store_cnt;
  wire   [5:0] out_cnt;
  wire   [2:0] out_cnt_6;
  wire   [1:0] m_size;
  wire   [5:0] in_cnt_64;
  wire   [7:0] in_cnt;
  wire   [3:0] in_matrix_cnt;
  wire   [63:0] in_64;
  wire   [9:0] in_addr_cnt;
  wire   [9:0] calin_addr;
  wire   [9:0] calweight_addr;
  wire   [3:0] i_mat;
  wire   [3:0] w_mat;
  wire   [8:0] in_start_addr;
  wire   [8:0] weight_start_addr;
  wire   [767:0] x_matrix;
  wire   [1023:0] w_matrix;
  wire   [7:0] cal_cnt;
  wire   [15:0] inA11;
  wire   [15:0] inA21;
  wire   [15:0] inA31;
  wire   [15:0] inA41;
  wire   [15:0] inA51;
  wire   [15:0] inA61;
  wire   [15:0] inA71;
  wire   [15:0] inA81;
  wire   [39:0] outC11;
  wire   [15:0] outD11;
  wire   [39:0] outC12;
  wire   [15:0] outD12;
  wire   [39:0] outC13;
  wire   [15:0] outD13;
  wire   [39:0] outC14;
  wire   [15:0] outD14;
  wire   [39:0] outC15;
  wire   [15:0] outD15;
  wire   [39:0] outC16;
  wire   [15:0] outD16;
  wire   [39:0] outC17;
  wire   [15:0] outD17;
  wire   [39:0] outC18;
  wire   [39:0] outC21;
  wire   [15:0] outD21;
  wire   [39:0] outC22;
  wire   [15:0] outD22;
  wire   [39:0] outC23;
  wire   [15:0] outD23;
  wire   [39:0] outC24;
  wire   [15:0] outD24;
  wire   [39:0] outC25;
  wire   [15:0] outD25;
  wire   [39:0] outC26;
  wire   [15:0] outD26;
  wire   [39:0] outC27;
  wire   [15:0] outD27;
  wire   [39:0] outC28;
  wire   [39:0] outC31;
  wire   [15:0] outD31;
  wire   [39:0] outC32;
  wire   [15:0] outD32;
  wire   [39:0] outC33;
  wire   [15:0] outD33;
  wire   [39:0] outC34;
  wire   [15:0] outD34;
  wire   [39:0] outC35;
  wire   [15:0] outD35;
  wire   [39:0] outC36;
  wire   [15:0] outD36;
  wire   [39:0] outC37;
  wire   [15:0] outD37;
  wire   [39:0] outC38;
  wire   [39:0] outC41;
  wire   [15:0] outD41;
  wire   [39:0] outC42;
  wire   [15:0] outD42;
  wire   [39:0] outC43;
  wire   [15:0] outD43;
  wire   [39:0] outC44;
  wire   [15:0] outD44;
  wire   [39:0] outC45;
  wire   [15:0] outD45;
  wire   [39:0] outC46;
  wire   [15:0] outD46;
  wire   [39:0] outC47;
  wire   [15:0] outD47;
  wire   [39:0] outC48;
  wire   [39:0] outC51;
  wire   [15:0] outD51;
  wire   [39:0] outC52;
  wire   [15:0] outD52;
  wire   [39:0] outC53;
  wire   [15:0] outD53;
  wire   [39:0] outC54;
  wire   [15:0] outD54;
  wire   [39:0] outC55;
  wire   [15:0] outD55;
  wire   [39:0] outC56;
  wire   [15:0] outD56;
  wire   [39:0] outC57;
  wire   [15:0] outD57;
  wire   [39:0] outC58;
  wire   [39:0] outC61;
  wire   [15:0] outD61;
  wire   [39:0] outC62;
  wire   [15:0] outD62;
  wire   [39:0] outC63;
  wire   [15:0] outD63;
  wire   [39:0] outC64;
  wire   [15:0] outD64;
  wire   [39:0] outC65;
  wire   [15:0] outD65;
  wire   [39:0] outC66;
  wire   [15:0] outD66;
  wire   [39:0] outC67;
  wire   [15:0] outD67;
  wire   [39:0] outC68;
  wire   [39:0] outC71;
  wire   [15:0] outD71;
  wire   [39:0] outC72;
  wire   [15:0] outD72;
  wire   [39:0] outC73;
  wire   [15:0] outD73;
  wire   [39:0] outC74;
  wire   [15:0] outD74;
  wire   [39:0] outC75;
  wire   [15:0] outD75;
  wire   [39:0] outC76;
  wire   [15:0] outD76;
  wire   [39:0] outC77;
  wire   [15:0] outD77;
  wire   [39:0] outC78;
  wire   [39:0] outC81;
  wire   [15:0] outD81;
  wire   [39:0] outC82;
  wire   [15:0] outD82;
  wire   [39:0] outC83;
  wire   [15:0] outD83;
  wire   [39:0] outC84;
  wire   [15:0] outD84;
  wire   [39:0] outC85;
  wire   [15:0] outD85;
  wire   [39:0] outC86;
  wire   [15:0] outD86;
  wire   [39:0] outC87;
  wire   [15:0] outD87;
  wire   [39:0] outC88;
  wire   [39:0] c_plus;
  wire   [599:0] cal_out;
  wire   [89:0] length_reg;
  wire   [39:0] value_out;
  wire   [5:0] length_out;
  wire   [4:2] add_250_carry;
  wire   [5:2] add_220_carry;
  tri   [63:0] mem_in_Q;
  tri   [63:0] mem_weight_Q;

  RA1SH MEM_IN ( .Q(mem_in_Q), .A({n5869, n5870, n5871, n5872, n5873, n5874, 
        n5875, n5876}), .D(in_64), .CLK(clk), .CEN(1'b0), .OEN(1'b0), .WEN(
        wen_in) );
  RA1SH MEM_WEIGHT ( .Q(mem_weight_Q), .A({n5861, n5862, n5863, n5864, n5865, 
        n5866, n5867, n5868}), .D(in_64), .CLK(clk), .CEN(1'b0), .OEN(1'b0), 
        .WEN(wen_weight) );
  NAND4X4 U2969 ( .A(n5821), .B(n5822), .C(n5823), .D(n754), .Y(n925) );
  OAI221X4 U3151 ( .A0(in_valid), .A1(n5066), .B0(n873), .B1(n1038), .C0(n1114), .Y(ns[2]) );
  AOI221X4 U3930 ( .A0(n1318), .A1(x_matrix[253]), .B0(n1384), .B1(
        x_matrix[349]), .C0(n1665), .Y(n1664) );
  AOI31X4 U3939 ( .A0(n1670), .A1(n1671), .A2(n1672), .B0(n1656), .Y(N11405)
         );
  AOI221X4 U3940 ( .A0(n1318), .A1(x_matrix[251]), .B0(n1384), .B1(
        x_matrix[347]), .C0(n1673), .Y(n1672) );
  AOI31X4 U3949 ( .A0(n1678), .A1(n1679), .A2(n1680), .B0(n1656), .Y(N11403)
         );
  AOI221X4 U3950 ( .A0(n1318), .A1(x_matrix[249]), .B0(n1384), .B1(
        x_matrix[345]), .C0(n1681), .Y(n1680) );
  AOI221X4 U3955 ( .A0(n1318), .A1(x_matrix[248]), .B0(n1384), .B1(
        x_matrix[344]), .C0(n1685), .Y(n1684) );
  AOI31X4 U3959 ( .A0(n1686), .A1(n1687), .A2(n1688), .B0(n1656), .Y(N11401)
         );
  AOI221X4 U3960 ( .A0(n1318), .A1(x_matrix[247]), .B0(n1384), .B1(
        x_matrix[343]), .C0(n1689), .Y(n1688) );
  AOI31X4 U3964 ( .A0(n1690), .A1(n1691), .A2(n1692), .B0(n1656), .Y(N11400)
         );
  AOI221X4 U3965 ( .A0(n1318), .A1(x_matrix[246]), .B0(n1384), .B1(
        x_matrix[342]), .C0(n1693), .Y(n1692) );
  AOI31X4 U3969 ( .A0(n1694), .A1(n1695), .A2(n1696), .B0(n1656), .Y(N11399)
         );
  AOI221X4 U3970 ( .A0(n1318), .A1(x_matrix[245]), .B0(n1384), .B1(
        x_matrix[341]), .C0(n1697), .Y(n1696) );
  AOI31X4 U3974 ( .A0(n1698), .A1(n1699), .A2(n1700), .B0(n1656), .Y(N11398)
         );
  AOI221X4 U3975 ( .A0(n1318), .A1(x_matrix[244]), .B0(n1384), .B1(
        x_matrix[340]), .C0(n1701), .Y(n1700) );
  AOI31X4 U3979 ( .A0(n1702), .A1(n1703), .A2(n1704), .B0(n1656), .Y(N11397)
         );
  AOI221X4 U3980 ( .A0(n1318), .A1(x_matrix[243]), .B0(n1384), .B1(
        x_matrix[339]), .C0(n1705), .Y(n1704) );
  AOI31X4 U3984 ( .A0(n1706), .A1(n1707), .A2(n1708), .B0(n1656), .Y(N11396)
         );
  AOI221X4 U3985 ( .A0(n1318), .A1(x_matrix[242]), .B0(n1384), .B1(
        x_matrix[338]), .C0(n1709), .Y(n1708) );
  AOI31X4 U3989 ( .A0(n1710), .A1(n1711), .A2(n1712), .B0(n1656), .Y(N11395)
         );
  AOI221X4 U3990 ( .A0(n1318), .A1(x_matrix[241]), .B0(n1384), .B1(
        x_matrix[337]), .C0(n1713), .Y(n1712) );
  AOI31X4 U3994 ( .A0(n1714), .A1(n1715), .A2(n1716), .B0(n1656), .Y(N11394)
         );
  AOI221X4 U3997 ( .A0(n1318), .A1(x_matrix[240]), .B0(n1384), .B1(
        x_matrix[336]), .C0(n1717), .Y(n1716) );
  NOR3X4 U4001 ( .A(cal_cnt[0]), .B(n5088), .C(n5893), .Y(n1384) );
  NOR3X4 U4002 ( .A(n5893), .B(n5088), .C(n5891), .Y(n1318) );
  PE_0 PE1_1 ( .rst_n(rst_n), .clk(clk), .inA(inA11), .inB({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .inW(w_matrix[1023:1008]), .outC(outC11), .outD(outD11) );
  PE_63 PE1_2 ( .rst_n(rst_n), .clk(clk), .inA(outD11), .inB({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .inW(w_matrix[1007:992]), .outC(outC12), .outD(outD12) );
  PE_62 PE1_3 ( .rst_n(rst_n), .clk(clk), .inA(outD12), .inB({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .inW(w_matrix[991:976]), .outC(outC13), .outD(outD13) );
  PE_61 PE1_4 ( .rst_n(rst_n), .clk(clk), .inA(outD13), .inB({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .inW(w_matrix[975:960]), .outC(outC14), .outD(outD14) );
  PE_60 PE1_5 ( .rst_n(rst_n), .clk(clk), .inA(outD14), .inB({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .inW(w_matrix[959:944]), .outC(outC15), .outD(outD15) );
  PE_59 PE1_6 ( .rst_n(rst_n), .clk(clk), .inA(outD15), .inB({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .inW(w_matrix[943:928]), .outC(outC16), .outD(outD16) );
  PE_58 PE1_7 ( .rst_n(rst_n), .clk(clk), .inA(outD16), .inB({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .inW(w_matrix[927:912]), .outC(outC17), .outD(outD17) );
  PE_57 PE1_8 ( .rst_n(rst_n), .clk(clk), .inA(outD17), .inB({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .inW(w_matrix[911:896]), .outC(outC18), .outD({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16}) );
  PE_56 PE2_1 ( .rst_n(rst_n), .clk(clk), .inA(inA21), .inB(outC11), .inW(
        w_matrix[895:880]), .outC(outC21), .outD(outD21) );
  PE_55 PE2_2 ( .rst_n(rst_n), .clk(clk), .inA(outD21), .inB(outC12), .inW(
        w_matrix[879:864]), .outC(outC22), .outD(outD22) );
  PE_54 PE2_3 ( .rst_n(rst_n), .clk(clk), .inA(outD22), .inB(outC13), .inW(
        w_matrix[863:848]), .outC(outC23), .outD(outD23) );
  PE_53 PE2_4 ( .rst_n(rst_n), .clk(clk), .inA(outD23), .inB(outC14), .inW(
        w_matrix[847:832]), .outC(outC24), .outD(outD24) );
  PE_52 PE2_5 ( .rst_n(rst_n), .clk(clk), .inA(outD24), .inB(outC15), .inW(
        w_matrix[831:816]), .outC(outC25), .outD(outD25) );
  PE_51 PE2_6 ( .rst_n(rst_n), .clk(clk), .inA(outD25), .inB(outC16), .inW(
        w_matrix[815:800]), .outC(outC26), .outD(outD26) );
  PE_50 PE2_7 ( .rst_n(rst_n), .clk(clk), .inA(outD26), .inB(outC17), .inW(
        w_matrix[799:784]), .outC(outC27), .outD(outD27) );
  PE_49 PE2_8 ( .rst_n(rst_n), .clk(clk), .inA(outD27), .inB(outC18), .inW(
        w_matrix[783:768]), .outC(outC28), .outD({SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32}) );
  PE_48 PE3_1 ( .rst_n(rst_n), .clk(clk), .inA(inA31), .inB(outC21), .inW(
        w_matrix[767:752]), .outC(outC31), .outD(outD31) );
  PE_47 PE3_2 ( .rst_n(rst_n), .clk(clk), .inA(outD31), .inB(outC22), .inW(
        w_matrix[751:736]), .outC(outC32), .outD(outD32) );
  PE_46 PE3_3 ( .rst_n(rst_n), .clk(clk), .inA(outD32), .inB(outC23), .inW(
        w_matrix[735:720]), .outC(outC33), .outD(outD33) );
  PE_45 PE3_4 ( .rst_n(rst_n), .clk(clk), .inA(outD33), .inB(outC24), .inW(
        w_matrix[719:704]), .outC(outC34), .outD(outD34) );
  PE_44 PE3_5 ( .rst_n(rst_n), .clk(clk), .inA(outD34), .inB(outC25), .inW(
        w_matrix[703:688]), .outC(outC35), .outD(outD35) );
  PE_43 PE3_6 ( .rst_n(rst_n), .clk(clk), .inA(outD35), .inB(outC26), .inW(
        w_matrix[687:672]), .outC(outC36), .outD(outD36) );
  PE_42 PE3_7 ( .rst_n(rst_n), .clk(clk), .inA(outD36), .inB(outC27), .inW(
        w_matrix[671:656]), .outC(outC37), .outD(outD37) );
  PE_41 PE3_8 ( .rst_n(rst_n), .clk(clk), .inA(outD37), .inB(outC28), .inW(
        w_matrix[655:640]), .outC(outC38), .outD({SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48}) );
  PE_40 PE4_1 ( .rst_n(rst_n), .clk(clk), .inA(inA41), .inB(outC31), .inW(
        w_matrix[639:624]), .outC(outC41), .outD(outD41) );
  PE_39 PE4_2 ( .rst_n(rst_n), .clk(clk), .inA(outD41), .inB(outC32), .inW(
        w_matrix[623:608]), .outC(outC42), .outD(outD42) );
  PE_38 PE4_3 ( .rst_n(rst_n), .clk(clk), .inA(outD42), .inB(outC33), .inW(
        w_matrix[607:592]), .outC(outC43), .outD(outD43) );
  PE_37 PE4_4 ( .rst_n(rst_n), .clk(clk), .inA(outD43), .inB(outC34), .inW(
        w_matrix[591:576]), .outC(outC44), .outD(outD44) );
  PE_36 PE4_5 ( .rst_n(rst_n), .clk(clk), .inA(outD44), .inB(outC35), .inW(
        w_matrix[575:560]), .outC(outC45), .outD(outD45) );
  PE_35 PE4_6 ( .rst_n(rst_n), .clk(clk), .inA(outD45), .inB(outC36), .inW(
        w_matrix[559:544]), .outC(outC46), .outD(outD46) );
  PE_34 PE4_7 ( .rst_n(rst_n), .clk(clk), .inA(outD46), .inB(outC37), .inW(
        w_matrix[543:528]), .outC(outC47), .outD(outD47) );
  PE_33 PE4_8 ( .rst_n(rst_n), .clk(clk), .inA(outD47), .inB(outC38), .inW(
        w_matrix[527:512]), .outC(outC48), .outD({SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64}) );
  PE_32 PE5_1 ( .rst_n(rst_n), .clk(clk), .inA(inA51), .inB(outC41), .inW(
        w_matrix[511:496]), .outC(outC51), .outD(outD51) );
  PE_31 PE5_2 ( .rst_n(rst_n), .clk(clk), .inA(outD51), .inB(outC42), .inW(
        w_matrix[495:480]), .outC(outC52), .outD(outD52) );
  PE_30 PE5_3 ( .rst_n(rst_n), .clk(clk), .inA(outD52), .inB(outC43), .inW(
        w_matrix[479:464]), .outC(outC53), .outD(outD53) );
  PE_29 PE5_4 ( .rst_n(rst_n), .clk(clk), .inA(outD53), .inB(outC44), .inW(
        w_matrix[463:448]), .outC(outC54), .outD(outD54) );
  PE_28 PE5_5 ( .rst_n(rst_n), .clk(clk), .inA(outD54), .inB(outC45), .inW(
        w_matrix[447:432]), .outC(outC55), .outD(outD55) );
  PE_27 PE5_6 ( .rst_n(rst_n), .clk(clk), .inA(outD55), .inB(outC46), .inW(
        w_matrix[431:416]), .outC(outC56), .outD(outD56) );
  PE_26 PE5_7 ( .rst_n(rst_n), .clk(clk), .inA(outD56), .inB(outC47), .inW(
        w_matrix[415:400]), .outC(outC57), .outD(outD57) );
  PE_25 PE5_8 ( .rst_n(rst_n), .clk(clk), .inA(outD57), .inB(outC48), .inW(
        w_matrix[399:384]), .outC(outC58), .outD({SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80}) );
  PE_24 PE6_1 ( .rst_n(rst_n), .clk(clk), .inA(inA61), .inB(outC51), .inW(
        w_matrix[383:368]), .outC(outC61), .outD(outD61) );
  PE_23 PE6_2 ( .rst_n(rst_n), .clk(clk), .inA(outD61), .inB(outC52), .inW(
        w_matrix[367:352]), .outC(outC62), .outD(outD62) );
  PE_22 PE6_3 ( .rst_n(rst_n), .clk(clk), .inA(outD62), .inB(outC53), .inW(
        w_matrix[351:336]), .outC(outC63), .outD(outD63) );
  PE_21 PE6_4 ( .rst_n(rst_n), .clk(clk), .inA(outD63), .inB(outC54), .inW(
        w_matrix[335:320]), .outC(outC64), .outD(outD64) );
  PE_20 PE6_5 ( .rst_n(rst_n), .clk(clk), .inA(outD64), .inB(outC55), .inW(
        w_matrix[319:304]), .outC(outC65), .outD(outD65) );
  PE_19 PE6_6 ( .rst_n(rst_n), .clk(clk), .inA(outD65), .inB(outC56), .inW(
        w_matrix[303:288]), .outC(outC66), .outD(outD66) );
  PE_18 PE6_7 ( .rst_n(rst_n), .clk(clk), .inA(outD66), .inB(outC57), .inW(
        w_matrix[287:272]), .outC(outC67), .outD(outD67) );
  PE_17 PE6_8 ( .rst_n(rst_n), .clk(clk), .inA(outD67), .inB(outC58), .inW(
        w_matrix[271:256]), .outC(outC68), .outD({SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96}) );
  PE_16 PE7_1 ( .rst_n(rst_n), .clk(clk), .inA(inA71), .inB(outC61), .inW(
        w_matrix[255:240]), .outC(outC71), .outD(outD71) );
  PE_15 PE7_2 ( .rst_n(rst_n), .clk(clk), .inA(outD71), .inB(outC62), .inW(
        w_matrix[239:224]), .outC(outC72), .outD(outD72) );
  PE_14 PE7_3 ( .rst_n(rst_n), .clk(clk), .inA(outD72), .inB(outC63), .inW(
        w_matrix[223:208]), .outC(outC73), .outD(outD73) );
  PE_13 PE7_4 ( .rst_n(rst_n), .clk(clk), .inA(outD73), .inB(outC64), .inW(
        w_matrix[207:192]), .outC(outC74), .outD(outD74) );
  PE_12 PE7_5 ( .rst_n(rst_n), .clk(clk), .inA(outD74), .inB(outC65), .inW(
        w_matrix[191:176]), .outC(outC75), .outD(outD75) );
  PE_11 PE7_6 ( .rst_n(rst_n), .clk(clk), .inA(outD75), .inB(outC66), .inW(
        w_matrix[175:160]), .outC(outC76), .outD(outD76) );
  PE_10 PE7_7 ( .rst_n(rst_n), .clk(clk), .inA(outD76), .inB(outC67), .inW(
        w_matrix[159:144]), .outC(outC77), .outD(outD77) );
  PE_9 PE7_8 ( .rst_n(rst_n), .clk(clk), .inA(outD77), .inB(outC68), .inW(
        w_matrix[143:128]), .outC(outC78), .outD({SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112}) );
  PE_8 PE8_1 ( .rst_n(rst_n), .clk(clk), .inA(inA81), .inB(outC71), .inW(
        w_matrix[127:112]), .outC(outC81), .outD(outD81) );
  PE_7 PE8_2 ( .rst_n(rst_n), .clk(clk), .inA(outD81), .inB(outC72), .inW(
        w_matrix[111:96]), .outC(outC82), .outD(outD82) );
  PE_6 PE8_3 ( .rst_n(rst_n), .clk(clk), .inA(outD82), .inB(outC73), .inW(
        w_matrix[95:80]), .outC(outC83), .outD(outD83) );
  PE_5 PE8_4 ( .rst_n(rst_n), .clk(clk), .inA(outD83), .inB(outC74), .inW(
        w_matrix[79:64]), .outC(outC84), .outD(outD84) );
  PE_4 PE8_5 ( .rst_n(rst_n), .clk(clk), .inA(outD84), .inB(outC75), .inW(
        w_matrix[63:48]), .outC(outC85), .outD(outD85) );
  PE_3 PE8_6 ( .rst_n(rst_n), .clk(clk), .inA(outD85), .inB(outC76), .inW(
        w_matrix[47:32]), .outC(outC86), .outD(outD86) );
  PE_2 PE8_7 ( .rst_n(rst_n), .clk(clk), .inA(outD86), .inB(outC77), .inW(
        w_matrix[31:16]), .outC(outC87), .outD(outD87) );
  PE_1 PE8_8 ( .rst_n(rst_n), .clk(clk), .inA(outD87), .inB(outC78), .inW(
        w_matrix[15:0]), .outC(outC88), .outD({SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128}) );
  MMSA_DW01_add_0 add_733 ( .A(outC21), .B(outC22), .CI(1'b0), .SUM({N12125, 
        N12124, N12123, N12122, N12121, N12120, N12119, N12118, N12117, N12116, 
        N12115, N12114, N12113, N12112, N12111, N12110, N12109, N12108, N12107, 
        N12106, N12105, N12104, N12103, N12102, N12101, N12100, N12099, N12098, 
        N12097, N12096, N12095, N12094, N12093, N12092, N12091, N12090, N12089, 
        N12088, N12087, N12086}) );
  MMSA_DW01_inc_0 add_463 ( .A({cal_cnt[7:4], n5086, n5087, n5088, cal_cnt[0]}), .SUM({N11313, N11312, N11311, N11310, N11309, N11308, N11307, N11306}) );
  MMSA_DW01_inc_1 add_384 ( .A(calin_cnt), .SUM({N1361, N1360, N1359, N1358, 
        N1357, N1356, N1355, N1354}) );
  MMSA_DW01_inc_2 add_372 ( .A(calweight_addr), .SUM({N1339, N1338, N1337, 
        N1336, N1335, N1334, N1333, N1332, N1331, N1330}) );
  MMSA_DW01_inc_3 add_357 ( .A(calin_addr), .SUM({N1311, N1310, N1309, N1308, 
        N1307, N1306, N1305, N1304, N1303, N1302}) );
  MMSA_DW01_inc_4 add_280 ( .A(in_addr_cnt), .SUM({N1252, N1251, N1250, N1249, 
        N1248, N1247, N1246, N1245, N1244, N1243}) );
  MMSA_DW01_inc_6 add_237 ( .A(in_cnt), .SUM({N1060, N1059, N1058, N1057, 
        N1056, N1055, N1054, N1053}) );
  MMSA_DW01_add_7 add_6_root_add_0_root_add_735_7 ( .A(outC81), .B(outC85), 
        .CI(1'b0), .SUM({N12405, N12404, N12403, N12402, N12401, N12400, 
        N12399, N12398, N12397, N12396, N12395, N12394, N12393, N12392, N12391, 
        N12390, N12389, N12388, N12387, N12386, N12385, N12384, N12383, N12382, 
        N12381, N12380, N12379, N12378, N12377, N12376, N12375, N12374, N12373, 
        N12372, N12371, N12370, N12369, N12368, N12367, N12366}) );
  MMSA_DW01_add_6 add_3_root_add_0_root_add_735_7 ( .A(outC86), .B(outC88), 
        .CI(1'b0), .SUM({N12325, N12324, N12323, N12322, N12321, N12320, 
        N12319, N12318, N12317, N12316, N12315, N12314, N12313, N12312, N12311, 
        N12310, N12309, N12308, N12307, N12306, N12305, N12304, N12303, N12302, 
        N12301, N12300, N12299, N12298, N12297, N12296, N12295, N12294, N12293, 
        N12292, N12291, N12290, N12289, N12288, N12287, N12286}) );
  MMSA_DW01_add_5 add_2_root_add_0_root_add_735_7 ( .A({N12405, N12404, N12403, 
        N12402, N12401, N12400, N12399, N12398, N12397, N12396, N12395, N12394, 
        N12393, N12392, N12391, N12390, N12389, N12388, N12387, N12386, N12385, 
        N12384, N12383, N12382, N12381, N12380, N12379, N12378, N12377, N12376, 
        N12375, N12374, N12373, N12372, N12371, N12370, N12369, N12368, N12367, 
        N12366}), .B({N12325, N12324, N12323, N12322, N12321, N12320, N12319, 
        N12318, N12317, N12316, N12315, N12314, N12313, N12312, N12311, N12310, 
        N12309, N12308, N12307, N12306, N12305, N12304, N12303, N12302, N12301, 
        N12300, N12299, N12298, N12297, N12296, N12295, N12294, N12293, N12292, 
        N12291, N12290, N12289, N12288, N12287, N12286}), .CI(1'b0), .SUM({
        N12285, N12284, N12283, N12282, N12281, N12280, N12279, N12278, N12277, 
        N12276, N12275, N12274, N12273, N12272, N12271, N12270, N12269, N12268, 
        N12267, N12266, N12265, N12264, N12263, N12262, N12261, N12260, N12259, 
        N12258, N12257, N12256, N12255, N12254, N12253, N12252, N12251, N12250, 
        N12249, N12248, N12247, N12246}) );
  MMSA_DW01_add_4 add_4_root_add_0_root_add_735_7 ( .A(outC82), .B(outC84), 
        .CI(1'b0), .SUM({N12485, N12484, N12483, N12482, N12481, N12480, 
        N12479, N12478, N12477, N12476, N12475, N12474, N12473, N12472, N12471, 
        N12470, N12469, N12468, N12467, N12466, N12465, N12464, N12463, N12462, 
        N12461, N12460, N12459, N12458, N12457, N12456, N12455, N12454, N12453, 
        N12452, N12451, N12450, N12449, N12448, N12447, N12446}) );
  MMSA_DW01_add_3 add_5_root_add_0_root_add_735_7 ( .A(outC83), .B(outC87), 
        .CI(1'b0), .SUM({N12365, N12364, N12363, N12362, N12361, N12360, 
        N12359, N12358, N12357, N12356, N12355, N12354, N12353, N12352, N12351, 
        N12350, N12349, N12348, N12347, N12346, N12345, N12344, N12343, N12342, 
        N12341, N12340, N12339, N12338, N12337, N12336, N12335, N12334, N12333, 
        N12332, N12331, N12330, N12329, N12328, N12327, N12326}) );
  MMSA_DW01_add_2 add_1_root_add_0_root_add_735_7 ( .A({N12485, N12484, N12483, 
        N12482, N12481, N12480, N12479, N12478, N12477, N12476, N12475, N12474, 
        N12473, N12472, N12471, N12470, N12469, N12468, N12467, N12466, N12465, 
        N12464, N12463, N12462, N12461, N12460, N12459, N12458, N12457, N12456, 
        N12455, N12454, N12453, N12452, N12451, N12450, N12449, N12448, N12447, 
        N12446}), .B({N12365, N12364, N12363, N12362, N12361, N12360, N12359, 
        N12358, N12357, N12356, N12355, N12354, N12353, N12352, N12351, N12350, 
        N12349, N12348, N12347, N12346, N12345, N12344, N12343, N12342, N12341, 
        N12340, N12339, N12338, N12337, N12336, N12335, N12334, N12333, N12332, 
        N12331, N12330, N12329, N12328, N12327, N12326}), .CI(1'b0), .SUM({
        N12445, N12444, N12443, N12442, N12441, N12440, N12439, N12438, N12437, 
        N12436, N12435, N12434, N12433, N12432, N12431, N12430, N12429, N12428, 
        N12427, N12426, N12425, N12424, N12423, N12422, N12421, N12420, N12419, 
        N12418, N12417, N12416, N12415, N12414, N12413, N12412, N12411, N12410, 
        N12409, N12408, N12407, N12406}) );
  MMSA_DW01_add_1 add_0_root_add_0_root_add_735_7 ( .A({N12285, N12284, N12283, 
        N12282, N12281, N12280, N12279, N12278, N12277, N12276, N12275, N12274, 
        N12273, N12272, N12271, N12270, N12269, N12268, N12267, N12266, N12265, 
        N12264, N12263, N12262, N12261, N12260, N12259, N12258, N12257, N12256, 
        N12255, N12254, N12253, N12252, N12251, N12250, N12249, N12248, N12247, 
        N12246}), .B({N12445, N12444, N12443, N12442, N12441, N12440, N12439, 
        N12438, N12437, N12436, N12435, N12434, N12433, N12432, N12431, N12430, 
        N12429, N12428, N12427, N12426, N12425, N12424, N12423, N12422, N12421, 
        N12420, N12419, N12418, N12417, N12416, N12415, N12414, N12413, N12412, 
        N12411, N12410, N12409, N12408, N12407, N12406}), .CI(1'b0), .SUM({
        N12525, N12524, N12523, N12522, N12521, N12520, N12519, N12518, N12517, 
        N12516, N12515, N12514, N12513, N12512, N12511, N12510, N12509, N12508, 
        N12507, N12506, N12505, N12504, N12503, N12502, N12501, N12500, N12499, 
        N12498, N12497, N12496, N12495, N12494, N12493, N12492, N12491, N12490, 
        N12489, N12488, N12487, N12486}) );
  MMSA_DW01_add_10 add_2_root_add_0_root_add_734_3 ( .A(outC41), .B(outC43), 
        .CI(1'b0), .SUM({N12205, N12204, N12203, N12202, N12201, N12200, 
        N12199, N12198, N12197, N12196, N12195, N12194, N12193, N12192, N12191, 
        N12190, N12189, N12188, N12187, N12186, N12185, N12184, N12183, N12182, 
        N12181, N12180, N12179, N12178, N12177, N12176, N12175, N12174, N12173, 
        N12172, N12171, N12170, N12169, N12168, N12167, N12166}) );
  MMSA_DW01_add_9 add_1_root_add_0_root_add_734_3 ( .A(outC42), .B(outC44), 
        .CI(1'b0), .SUM({N12165, N12164, N12163, N12162, N12161, N12160, 
        N12159, N12158, N12157, N12156, N12155, N12154, N12153, N12152, N12151, 
        N12150, N12149, N12148, N12147, N12146, N12145, N12144, N12143, N12142, 
        N12141, N12140, N12139, N12138, N12137, N12136, N12135, N12134, N12133, 
        N12132, N12131, N12130, N12129, N12128, N12127, N12126}) );
  MMSA_DW01_add_8 add_0_root_add_0_root_add_734_3 ( .A({N12205, N12204, N12203, 
        N12202, N12201, N12200, N12199, N12198, N12197, N12196, N12195, N12194, 
        N12193, N12192, N12191, N12190, N12189, N12188, N12187, N12186, N12185, 
        N12184, N12183, N12182, N12181, N12180, N12179, N12178, N12177, N12176, 
        N12175, N12174, N12173, N12172, N12171, N12170, N12169, N12168, N12167, 
        N12166}), .B({N12165, N12164, N12163, N12162, N12161, N12160, N12159, 
        N12158, N12157, N12156, N12155, N12154, N12153, N12152, N12151, N12150, 
        N12149, N12148, N12147, N12146, N12145, N12144, N12143, N12142, N12141, 
        N12140, N12139, N12138, N12137, N12136, N12135, N12134, N12133, N12132, 
        N12131, N12130, N12129, N12128, N12127, N12126}), .CI(1'b0), .SUM({
        N12245, N12244, N12243, N12242, N12241, N12240, N12239, N12238, N12237, 
        N12236, N12235, N12234, N12233, N12232, N12231, N12230, N12229, N12228, 
        N12227, N12226, N12225, N12224, N12223, N12222, N12221, N12220, N12219, 
        N12218, N12217, N12216, N12215, N12214, N12213, N12212, N12211, N12210, 
        N12209, N12208, N12207, N12206}) );
  MMSA_DW_mult_uns_1 mult_343 ( .a(w_mat), .b({n5064, 1'b0, n5061, 1'b0, 
        mem_num_0}), .product(weight_start_addr) );
  MMSA_DW_mult_uns_0 mult_342 ( .a(i_mat), .b({n5064, 1'b0, n5061, 1'b0, 
        mem_num_0}), .product(in_start_addr) );
  DFFRHQX1 in_64_reg_0_ ( .D(N1162), .CK(clk), .RN(rst_n), .Q(in_64[0]) );
  DFFRHQX1 in_64_reg_1_ ( .D(N1163), .CK(clk), .RN(rst_n), .Q(in_64[1]) );
  DFFRHQX1 in_64_reg_2_ ( .D(N1164), .CK(clk), .RN(rst_n), .Q(in_64[2]) );
  DFFRHQX1 in_64_reg_3_ ( .D(N1165), .CK(clk), .RN(rst_n), .Q(in_64[3]) );
  DFFRHQX1 in_64_reg_4_ ( .D(N1166), .CK(clk), .RN(rst_n), .Q(in_64[4]) );
  DFFRHQX1 in_64_reg_5_ ( .D(N1167), .CK(clk), .RN(rst_n), .Q(in_64[5]) );
  DFFRHQX1 in_64_reg_6_ ( .D(N1168), .CK(clk), .RN(rst_n), .Q(in_64[6]) );
  DFFRHQX1 in_64_reg_7_ ( .D(N1169), .CK(clk), .RN(rst_n), .Q(in_64[7]) );
  DFFRHQX1 in_64_reg_8_ ( .D(N1170), .CK(clk), .RN(rst_n), .Q(in_64[8]) );
  DFFRHQX1 in_64_reg_9_ ( .D(N1171), .CK(clk), .RN(rst_n), .Q(in_64[9]) );
  DFFRHQX1 in_64_reg_10_ ( .D(N1172), .CK(clk), .RN(rst_n), .Q(in_64[10]) );
  DFFRHQX1 in_64_reg_11_ ( .D(N1173), .CK(clk), .RN(rst_n), .Q(in_64[11]) );
  DFFRHQX1 in_64_reg_12_ ( .D(N1174), .CK(clk), .RN(rst_n), .Q(in_64[12]) );
  DFFRHQX1 in_64_reg_13_ ( .D(N1175), .CK(clk), .RN(rst_n), .Q(in_64[13]) );
  DFFRHQX1 in_64_reg_14_ ( .D(N1176), .CK(clk), .RN(rst_n), .Q(in_64[14]) );
  DFFRHQX1 in_64_reg_15_ ( .D(N1177), .CK(clk), .RN(rst_n), .Q(in_64[15]) );
  DFFRHQX1 in_64_reg_16_ ( .D(N1178), .CK(clk), .RN(rst_n), .Q(in_64[16]) );
  DFFRHQX1 in_64_reg_17_ ( .D(N1179), .CK(clk), .RN(rst_n), .Q(in_64[17]) );
  DFFRHQX1 in_64_reg_18_ ( .D(N1180), .CK(clk), .RN(rst_n), .Q(in_64[18]) );
  DFFRHQX1 in_64_reg_19_ ( .D(N1181), .CK(clk), .RN(rst_n), .Q(in_64[19]) );
  DFFRHQX1 in_64_reg_20_ ( .D(N1182), .CK(clk), .RN(rst_n), .Q(in_64[20]) );
  DFFRHQX1 in_64_reg_21_ ( .D(N1183), .CK(clk), .RN(rst_n), .Q(in_64[21]) );
  DFFRHQX1 in_64_reg_22_ ( .D(N1184), .CK(clk), .RN(rst_n), .Q(in_64[22]) );
  DFFRHQX1 in_64_reg_23_ ( .D(N1185), .CK(clk), .RN(rst_n), .Q(in_64[23]) );
  DFFRHQX1 in_64_reg_24_ ( .D(N1186), .CK(clk), .RN(rst_n), .Q(in_64[24]) );
  DFFRHQX1 in_64_reg_25_ ( .D(N1187), .CK(clk), .RN(rst_n), .Q(in_64[25]) );
  DFFRHQX1 in_64_reg_26_ ( .D(N1188), .CK(clk), .RN(rst_n), .Q(in_64[26]) );
  DFFRHQX1 in_64_reg_27_ ( .D(N1189), .CK(clk), .RN(rst_n), .Q(in_64[27]) );
  DFFRHQX1 in_64_reg_28_ ( .D(N1190), .CK(clk), .RN(rst_n), .Q(in_64[28]) );
  DFFRHQX1 in_64_reg_29_ ( .D(N1191), .CK(clk), .RN(rst_n), .Q(in_64[29]) );
  DFFRHQX1 in_64_reg_30_ ( .D(N1192), .CK(clk), .RN(rst_n), .Q(in_64[30]) );
  DFFRHQX1 in_64_reg_31_ ( .D(N1193), .CK(clk), .RN(rst_n), .Q(in_64[31]) );
  DFFRHQX1 in_64_reg_32_ ( .D(N1194), .CK(clk), .RN(rst_n), .Q(in_64[32]) );
  DFFRHQX1 in_64_reg_33_ ( .D(N1195), .CK(clk), .RN(rst_n), .Q(in_64[33]) );
  DFFRHQX1 in_64_reg_34_ ( .D(N1196), .CK(clk), .RN(rst_n), .Q(in_64[34]) );
  DFFRHQX1 in_64_reg_35_ ( .D(N1197), .CK(clk), .RN(rst_n), .Q(in_64[35]) );
  DFFRHQX1 in_64_reg_36_ ( .D(N1198), .CK(clk), .RN(rst_n), .Q(in_64[36]) );
  DFFRHQX1 in_64_reg_37_ ( .D(N1199), .CK(clk), .RN(rst_n), .Q(in_64[37]) );
  DFFRHQX1 in_64_reg_38_ ( .D(N1200), .CK(clk), .RN(rst_n), .Q(in_64[38]) );
  DFFRHQX1 in_64_reg_39_ ( .D(N1201), .CK(clk), .RN(rst_n), .Q(in_64[39]) );
  DFFRHQX1 in_64_reg_40_ ( .D(N1202), .CK(clk), .RN(rst_n), .Q(in_64[40]) );
  DFFRHQX1 in_64_reg_41_ ( .D(N1203), .CK(clk), .RN(rst_n), .Q(in_64[41]) );
  DFFRHQX1 in_64_reg_42_ ( .D(N1204), .CK(clk), .RN(rst_n), .Q(in_64[42]) );
  DFFRHQX1 in_64_reg_43_ ( .D(N1205), .CK(clk), .RN(rst_n), .Q(in_64[43]) );
  DFFRHQX1 in_64_reg_44_ ( .D(N1206), .CK(clk), .RN(rst_n), .Q(in_64[44]) );
  DFFRHQX1 in_64_reg_45_ ( .D(N1207), .CK(clk), .RN(rst_n), .Q(in_64[45]) );
  DFFRHQX1 in_64_reg_46_ ( .D(N1208), .CK(clk), .RN(rst_n), .Q(in_64[46]) );
  DFFRHQX1 in_64_reg_47_ ( .D(N1209), .CK(clk), .RN(rst_n), .Q(in_64[47]) );
  DFFRHQX1 in_64_reg_48_ ( .D(N1210), .CK(clk), .RN(rst_n), .Q(in_64[48]) );
  DFFRHQX1 in_64_reg_49_ ( .D(N1211), .CK(clk), .RN(rst_n), .Q(in_64[49]) );
  DFFRHQX1 in_64_reg_50_ ( .D(N1212), .CK(clk), .RN(rst_n), .Q(in_64[50]) );
  DFFRHQX1 in_64_reg_51_ ( .D(N1213), .CK(clk), .RN(rst_n), .Q(in_64[51]) );
  DFFRHQX1 in_64_reg_52_ ( .D(N1214), .CK(clk), .RN(rst_n), .Q(in_64[52]) );
  DFFRHQX1 in_64_reg_53_ ( .D(N1215), .CK(clk), .RN(rst_n), .Q(in_64[53]) );
  DFFRHQX1 in_64_reg_54_ ( .D(N1216), .CK(clk), .RN(rst_n), .Q(in_64[54]) );
  DFFRHQX1 in_64_reg_55_ ( .D(N1217), .CK(clk), .RN(rst_n), .Q(in_64[55]) );
  DFFRHQX1 in_64_reg_56_ ( .D(N1218), .CK(clk), .RN(rst_n), .Q(in_64[56]) );
  DFFRHQX1 in_64_reg_57_ ( .D(N1219), .CK(clk), .RN(rst_n), .Q(in_64[57]) );
  DFFRHQX1 in_64_reg_58_ ( .D(N1220), .CK(clk), .RN(rst_n), .Q(in_64[58]) );
  DFFRHQX1 in_64_reg_59_ ( .D(N1221), .CK(clk), .RN(rst_n), .Q(in_64[59]) );
  DFFRHQX1 in_64_reg_60_ ( .D(N1222), .CK(clk), .RN(rst_n), .Q(in_64[60]) );
  DFFRHQX1 in_64_reg_61_ ( .D(N1223), .CK(clk), .RN(rst_n), .Q(in_64[61]) );
  DFFRHQX1 in_64_reg_62_ ( .D(N1224), .CK(clk), .RN(rst_n), .Q(in_64[62]) );
  DFFRHQX1 calweight_addr_reg_9_ ( .D(N1349), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[9]) );
  DFFRHQX1 calin_addr_reg_9_ ( .D(N1321), .CK(clk), .RN(rst_n), .Q(
        calin_addr[9]) );
  DFFRHQX1 x_matrix_reg_2__7__9_ ( .D(n3810), .CK(clk), .RN(rst_n), .Q(
        x_matrix[457]) );
  DFFRHQX1 x_matrix_reg_6__3__9_ ( .D(n4258), .CK(clk), .RN(rst_n), .Q(
        x_matrix[153]) );
  DFFRHQX1 x_matrix_reg_2__7__8_ ( .D(n3811), .CK(clk), .RN(rst_n), .Q(
        x_matrix[456]) );
  DFFRHQX1 x_matrix_reg_6__3__8_ ( .D(n4259), .CK(clk), .RN(rst_n), .Q(
        x_matrix[152]) );
  DFFRHQX1 x_matrix_reg_2__7__7_ ( .D(n3812), .CK(clk), .RN(rst_n), .Q(
        x_matrix[455]) );
  DFFRHQX1 x_matrix_reg_6__3__7_ ( .D(n4260), .CK(clk), .RN(rst_n), .Q(
        x_matrix[151]) );
  DFFRHQX1 x_matrix_reg_2__7__6_ ( .D(n3813), .CK(clk), .RN(rst_n), .Q(
        x_matrix[454]) );
  DFFRHQX1 x_matrix_reg_6__3__6_ ( .D(n4261), .CK(clk), .RN(rst_n), .Q(
        x_matrix[150]) );
  DFFRHQX1 x_matrix_reg_4__0__15_ ( .D(n3948), .CK(clk), .RN(rst_n), .Q(
        x_matrix[351]) );
  DFFRHQX1 x_matrix_reg_6__4__15_ ( .D(n4268), .CK(clk), .RN(rst_n), .Q(
        x_matrix[143]) );
  DFFRHQX1 x_matrix_reg_4__0__14_ ( .D(n3949), .CK(clk), .RN(rst_n), .Q(
        x_matrix[350]) );
  DFFRHQX1 x_matrix_reg_6__4__14_ ( .D(n4269), .CK(clk), .RN(rst_n), .Q(
        x_matrix[142]) );
  DFFRHQX1 x_matrix_reg_4__0__13_ ( .D(n3950), .CK(clk), .RN(rst_n), .Q(
        x_matrix[349]) );
  DFFRHQX1 x_matrix_reg_6__4__13_ ( .D(n4270), .CK(clk), .RN(rst_n), .Q(
        x_matrix[141]) );
  DFFRHQX1 x_matrix_reg_4__0__12_ ( .D(n3951), .CK(clk), .RN(rst_n), .Q(
        x_matrix[348]) );
  DFFRHQX1 x_matrix_reg_6__4__12_ ( .D(n4271), .CK(clk), .RN(rst_n), .Q(
        x_matrix[140]) );
  DFFRHQX1 x_matrix_reg_2__7__5_ ( .D(n3814), .CK(clk), .RN(rst_n), .Q(
        x_matrix[453]) );
  DFFRHQX1 x_matrix_reg_6__3__5_ ( .D(n4262), .CK(clk), .RN(rst_n), .Q(
        x_matrix[149]) );
  DFFRHQX1 x_matrix_reg_4__0__11_ ( .D(n3952), .CK(clk), .RN(rst_n), .Q(
        x_matrix[347]) );
  DFFRHQX1 x_matrix_reg_6__4__11_ ( .D(n4272), .CK(clk), .RN(rst_n), .Q(
        x_matrix[139]) );
  DFFRHQX1 x_matrix_reg_4__0__10_ ( .D(n3953), .CK(clk), .RN(rst_n), .Q(
        x_matrix[346]) );
  DFFRHQX1 x_matrix_reg_6__4__10_ ( .D(n4273), .CK(clk), .RN(rst_n), .Q(
        x_matrix[138]) );
  DFFRHQX1 x_matrix_reg_4__0__9_ ( .D(n3954), .CK(clk), .RN(rst_n), .Q(
        x_matrix[345]) );
  DFFRHQX1 x_matrix_reg_6__4__9_ ( .D(n4274), .CK(clk), .RN(rst_n), .Q(
        x_matrix[137]) );
  DFFRHQX1 x_matrix_reg_4__0__8_ ( .D(n3955), .CK(clk), .RN(rst_n), .Q(
        x_matrix[344]) );
  DFFRHQX1 x_matrix_reg_6__4__8_ ( .D(n4275), .CK(clk), .RN(rst_n), .Q(
        x_matrix[136]) );
  DFFRHQX1 x_matrix_reg_4__0__7_ ( .D(n3956), .CK(clk), .RN(rst_n), .Q(
        x_matrix[343]) );
  DFFRHQX1 x_matrix_reg_6__4__7_ ( .D(n4276), .CK(clk), .RN(rst_n), .Q(
        x_matrix[135]) );
  DFFRHQX1 x_matrix_reg_4__0__6_ ( .D(n3957), .CK(clk), .RN(rst_n), .Q(
        x_matrix[342]) );
  DFFRHQX1 x_matrix_reg_6__4__6_ ( .D(n4277), .CK(clk), .RN(rst_n), .Q(
        x_matrix[134]) );
  DFFRHQX1 x_matrix_reg_4__0__5_ ( .D(n3958), .CK(clk), .RN(rst_n), .Q(
        x_matrix[341]) );
  DFFRHQX1 x_matrix_reg_6__4__5_ ( .D(n4278), .CK(clk), .RN(rst_n), .Q(
        x_matrix[133]) );
  DFFRHQX1 x_matrix_reg_4__0__4_ ( .D(n3959), .CK(clk), .RN(rst_n), .Q(
        x_matrix[340]) );
  DFFRHQX1 x_matrix_reg_6__4__4_ ( .D(n4279), .CK(clk), .RN(rst_n), .Q(
        x_matrix[132]) );
  DFFRHQX1 x_matrix_reg_4__0__3_ ( .D(n3960), .CK(clk), .RN(rst_n), .Q(
        x_matrix[339]) );
  DFFRHQX1 x_matrix_reg_6__4__3_ ( .D(n4280), .CK(clk), .RN(rst_n), .Q(
        x_matrix[131]) );
  DFFRHQX1 x_matrix_reg_4__0__2_ ( .D(n3961), .CK(clk), .RN(rst_n), .Q(
        x_matrix[338]) );
  DFFRHQX1 x_matrix_reg_6__4__2_ ( .D(n4281), .CK(clk), .RN(rst_n), .Q(
        x_matrix[130]) );
  DFFRHQX1 x_matrix_reg_2__7__4_ ( .D(n3815), .CK(clk), .RN(rst_n), .Q(
        x_matrix[452]) );
  DFFRHQX1 x_matrix_reg_6__3__4_ ( .D(n4263), .CK(clk), .RN(rst_n), .Q(
        x_matrix[148]) );
  DFFRHQX1 x_matrix_reg_4__0__1_ ( .D(n3962), .CK(clk), .RN(rst_n), .Q(
        x_matrix[337]) );
  DFFRHQX1 x_matrix_reg_6__4__1_ ( .D(n4282), .CK(clk), .RN(rst_n), .Q(
        x_matrix[129]) );
  DFFRHQX1 x_matrix_reg_4__0__0_ ( .D(n3963), .CK(clk), .RN(rst_n), .Q(
        x_matrix[336]) );
  DFFRHQX1 x_matrix_reg_6__4__0_ ( .D(n4283), .CK(clk), .RN(rst_n), .Q(
        x_matrix[128]) );
  DFFRHQX1 x_matrix_reg_0__5__15_ ( .D(n3516), .CK(clk), .RN(rst_n), .Q(
        x_matrix[687]) );
  DFFRHQX1 x_matrix_reg_4__1__15_ ( .D(n3964), .CK(clk), .RN(rst_n), .Q(
        x_matrix[335]) );
  DFFRHQX1 x_matrix_reg_0__5__14_ ( .D(n3517), .CK(clk), .RN(rst_n), .Q(
        x_matrix[686]) );
  DFFRHQX1 x_matrix_reg_4__1__14_ ( .D(n3965), .CK(clk), .RN(rst_n), .Q(
        x_matrix[334]) );
  DFFRHQX1 x_matrix_reg_0__5__13_ ( .D(n3518), .CK(clk), .RN(rst_n), .Q(
        x_matrix[685]) );
  DFFRHQX1 x_matrix_reg_4__1__13_ ( .D(n3966), .CK(clk), .RN(rst_n), .Q(
        x_matrix[333]) );
  DFFRHQX1 x_matrix_reg_0__5__12_ ( .D(n3519), .CK(clk), .RN(rst_n), .Q(
        x_matrix[684]) );
  DFFRHQX1 x_matrix_reg_4__1__12_ ( .D(n3967), .CK(clk), .RN(rst_n), .Q(
        x_matrix[332]) );
  DFFRHQX1 x_matrix_reg_0__5__11_ ( .D(n3520), .CK(clk), .RN(rst_n), .Q(
        x_matrix[683]) );
  DFFRHQX1 x_matrix_reg_4__1__11_ ( .D(n3968), .CK(clk), .RN(rst_n), .Q(
        x_matrix[331]) );
  DFFRHQX1 x_matrix_reg_0__5__10_ ( .D(n3521), .CK(clk), .RN(rst_n), .Q(
        x_matrix[682]) );
  DFFRHQX1 x_matrix_reg_4__1__10_ ( .D(n3969), .CK(clk), .RN(rst_n), .Q(
        x_matrix[330]) );
  DFFRHQX1 x_matrix_reg_0__5__9_ ( .D(n3522), .CK(clk), .RN(rst_n), .Q(
        x_matrix[681]) );
  DFFRHQX1 x_matrix_reg_4__1__9_ ( .D(n3970), .CK(clk), .RN(rst_n), .Q(
        x_matrix[329]) );
  DFFRHQX1 x_matrix_reg_0__5__8_ ( .D(n3523), .CK(clk), .RN(rst_n), .Q(
        x_matrix[680]) );
  DFFRHQX1 x_matrix_reg_4__1__8_ ( .D(n3971), .CK(clk), .RN(rst_n), .Q(
        x_matrix[328]) );
  DFFRHQX1 x_matrix_reg_2__7__3_ ( .D(n3816), .CK(clk), .RN(rst_n), .Q(
        x_matrix[451]) );
  DFFRHQX1 x_matrix_reg_6__3__3_ ( .D(n4264), .CK(clk), .RN(rst_n), .Q(
        x_matrix[147]) );
  DFFRHQX1 x_matrix_reg_0__5__7_ ( .D(n3524), .CK(clk), .RN(rst_n), .Q(
        x_matrix[679]) );
  DFFRHQX1 x_matrix_reg_4__1__7_ ( .D(n3972), .CK(clk), .RN(rst_n), .Q(
        x_matrix[327]) );
  DFFRHQX1 x_matrix_reg_0__5__6_ ( .D(n3525), .CK(clk), .RN(rst_n), .Q(
        x_matrix[678]) );
  DFFRHQX1 x_matrix_reg_4__1__6_ ( .D(n3973), .CK(clk), .RN(rst_n), .Q(
        x_matrix[326]) );
  DFFRHQX1 x_matrix_reg_0__5__5_ ( .D(n3526), .CK(clk), .RN(rst_n), .Q(
        x_matrix[677]) );
  DFFRHQX1 x_matrix_reg_4__1__5_ ( .D(n3974), .CK(clk), .RN(rst_n), .Q(
        x_matrix[325]) );
  DFFRHQX1 x_matrix_reg_0__5__4_ ( .D(n3527), .CK(clk), .RN(rst_n), .Q(
        x_matrix[676]) );
  DFFRHQX1 x_matrix_reg_4__1__4_ ( .D(n3975), .CK(clk), .RN(rst_n), .Q(
        x_matrix[324]) );
  DFFRHQX1 x_matrix_reg_0__5__3_ ( .D(n3528), .CK(clk), .RN(rst_n), .Q(
        x_matrix[675]) );
  DFFRHQX1 x_matrix_reg_4__1__3_ ( .D(n3976), .CK(clk), .RN(rst_n), .Q(
        x_matrix[323]) );
  DFFRHQX1 x_matrix_reg_0__5__2_ ( .D(n3529), .CK(clk), .RN(rst_n), .Q(
        x_matrix[674]) );
  DFFRHQX1 x_matrix_reg_4__1__2_ ( .D(n3977), .CK(clk), .RN(rst_n), .Q(
        x_matrix[322]) );
  DFFRHQX1 x_matrix_reg_0__5__1_ ( .D(n3530), .CK(clk), .RN(rst_n), .Q(
        x_matrix[673]) );
  DFFRHQX1 x_matrix_reg_4__1__1_ ( .D(n3978), .CK(clk), .RN(rst_n), .Q(
        x_matrix[321]) );
  DFFRHQX1 x_matrix_reg_0__5__0_ ( .D(n3531), .CK(clk), .RN(rst_n), .Q(
        x_matrix[672]) );
  DFFRHQX1 x_matrix_reg_4__1__0_ ( .D(n3979), .CK(clk), .RN(rst_n), .Q(
        x_matrix[320]) );
  DFFRHQX1 x_matrix_reg_0__6__15_ ( .D(n3532), .CK(clk), .RN(rst_n), .Q(
        x_matrix[671]) );
  DFFRHQX1 x_matrix_reg_4__2__15_ ( .D(n3980), .CK(clk), .RN(rst_n), .Q(
        x_matrix[319]) );
  DFFRHQX1 x_matrix_reg_0__6__14_ ( .D(n3533), .CK(clk), .RN(rst_n), .Q(
        x_matrix[670]) );
  DFFRHQX1 x_matrix_reg_4__2__14_ ( .D(n3981), .CK(clk), .RN(rst_n), .Q(
        x_matrix[318]) );
  DFFRHQX1 x_matrix_reg_2__7__2_ ( .D(n3817), .CK(clk), .RN(rst_n), .Q(
        x_matrix[450]) );
  DFFRHQX1 x_matrix_reg_6__3__2_ ( .D(n4265), .CK(clk), .RN(rst_n), .Q(
        x_matrix[146]) );
  DFFRHQX1 x_matrix_reg_0__6__13_ ( .D(n3534), .CK(clk), .RN(rst_n), .Q(
        x_matrix[669]) );
  DFFRHQX1 x_matrix_reg_4__2__13_ ( .D(n3982), .CK(clk), .RN(rst_n), .Q(
        x_matrix[317]) );
  DFFRHQX1 x_matrix_reg_0__6__12_ ( .D(n3535), .CK(clk), .RN(rst_n), .Q(
        x_matrix[668]) );
  DFFRHQX1 x_matrix_reg_4__2__12_ ( .D(n3983), .CK(clk), .RN(rst_n), .Q(
        x_matrix[316]) );
  DFFRHQX1 x_matrix_reg_0__6__11_ ( .D(n3536), .CK(clk), .RN(rst_n), .Q(
        x_matrix[667]) );
  DFFRHQX1 x_matrix_reg_4__2__11_ ( .D(n3984), .CK(clk), .RN(rst_n), .Q(
        x_matrix[315]) );
  DFFRHQX1 x_matrix_reg_0__6__10_ ( .D(n3537), .CK(clk), .RN(rst_n), .Q(
        x_matrix[666]) );
  DFFRHQX1 x_matrix_reg_4__2__10_ ( .D(n3985), .CK(clk), .RN(rst_n), .Q(
        x_matrix[314]) );
  DFFRHQX1 x_matrix_reg_0__6__9_ ( .D(n3538), .CK(clk), .RN(rst_n), .Q(
        x_matrix[665]) );
  DFFRHQX1 x_matrix_reg_4__2__9_ ( .D(n3986), .CK(clk), .RN(rst_n), .Q(
        x_matrix[313]) );
  DFFRHQX1 x_matrix_reg_0__6__8_ ( .D(n3539), .CK(clk), .RN(rst_n), .Q(
        x_matrix[664]) );
  DFFRHQX1 x_matrix_reg_4__2__8_ ( .D(n3987), .CK(clk), .RN(rst_n), .Q(
        x_matrix[312]) );
  DFFRHQX1 x_matrix_reg_0__6__7_ ( .D(n3540), .CK(clk), .RN(rst_n), .Q(
        x_matrix[663]) );
  DFFRHQX1 x_matrix_reg_4__2__7_ ( .D(n3988), .CK(clk), .RN(rst_n), .Q(
        x_matrix[311]) );
  DFFRHQX1 x_matrix_reg_0__6__6_ ( .D(n3541), .CK(clk), .RN(rst_n), .Q(
        x_matrix[662]) );
  DFFRHQX1 x_matrix_reg_4__2__6_ ( .D(n3989), .CK(clk), .RN(rst_n), .Q(
        x_matrix[310]) );
  DFFRHQX1 x_matrix_reg_0__6__5_ ( .D(n3542), .CK(clk), .RN(rst_n), .Q(
        x_matrix[661]) );
  DFFRHQX1 x_matrix_reg_4__2__5_ ( .D(n3990), .CK(clk), .RN(rst_n), .Q(
        x_matrix[309]) );
  DFFRHQX1 x_matrix_reg_0__6__4_ ( .D(n3543), .CK(clk), .RN(rst_n), .Q(
        x_matrix[660]) );
  DFFRHQX1 x_matrix_reg_4__2__4_ ( .D(n3991), .CK(clk), .RN(rst_n), .Q(
        x_matrix[308]) );
  DFFRHQX1 x_matrix_reg_2__7__1_ ( .D(n3818), .CK(clk), .RN(rst_n), .Q(
        x_matrix[449]) );
  DFFRHQX1 x_matrix_reg_6__3__1_ ( .D(n4266), .CK(clk), .RN(rst_n), .Q(
        x_matrix[145]) );
  DFFRHQX1 x_matrix_reg_0__6__3_ ( .D(n3544), .CK(clk), .RN(rst_n), .Q(
        x_matrix[659]) );
  DFFRHQX1 x_matrix_reg_4__2__3_ ( .D(n3992), .CK(clk), .RN(rst_n), .Q(
        x_matrix[307]) );
  DFFRHQX1 x_matrix_reg_0__6__2_ ( .D(n3545), .CK(clk), .RN(rst_n), .Q(
        x_matrix[658]) );
  DFFRHQX1 x_matrix_reg_4__2__2_ ( .D(n3993), .CK(clk), .RN(rst_n), .Q(
        x_matrix[306]) );
  DFFRHQX1 x_matrix_reg_0__6__1_ ( .D(n3546), .CK(clk), .RN(rst_n), .Q(
        x_matrix[657]) );
  DFFRHQX1 x_matrix_reg_4__2__1_ ( .D(n3994), .CK(clk), .RN(rst_n), .Q(
        x_matrix[305]) );
  DFFRHQX1 x_matrix_reg_0__6__0_ ( .D(n3547), .CK(clk), .RN(rst_n), .Q(
        x_matrix[656]) );
  DFFRHQX1 x_matrix_reg_4__2__0_ ( .D(n3995), .CK(clk), .RN(rst_n), .Q(
        x_matrix[304]) );
  DFFRHQX1 x_matrix_reg_2__7__15_ ( .D(n3804), .CK(clk), .RN(rst_n), .Q(
        x_matrix[463]) );
  DFFRHQX1 x_matrix_reg_6__3__15_ ( .D(n4252), .CK(clk), .RN(rst_n), .Q(
        x_matrix[159]) );
  DFFRHQX1 x_matrix_reg_2__7__14_ ( .D(n3805), .CK(clk), .RN(rst_n), .Q(
        x_matrix[462]) );
  DFFRHQX1 x_matrix_reg_6__3__14_ ( .D(n4253), .CK(clk), .RN(rst_n), .Q(
        x_matrix[158]) );
  DFFRHQX1 x_matrix_reg_2__7__13_ ( .D(n3806), .CK(clk), .RN(rst_n), .Q(
        x_matrix[461]) );
  DFFRHQX1 x_matrix_reg_6__3__13_ ( .D(n4254), .CK(clk), .RN(rst_n), .Q(
        x_matrix[157]) );
  DFFRHQX1 x_matrix_reg_2__7__12_ ( .D(n3807), .CK(clk), .RN(rst_n), .Q(
        x_matrix[460]) );
  DFFRHQX1 x_matrix_reg_6__3__12_ ( .D(n4255), .CK(clk), .RN(rst_n), .Q(
        x_matrix[156]) );
  DFFRHQX1 x_matrix_reg_2__7__11_ ( .D(n3808), .CK(clk), .RN(rst_n), .Q(
        x_matrix[459]) );
  DFFRHQX1 x_matrix_reg_6__3__11_ ( .D(n4256), .CK(clk), .RN(rst_n), .Q(
        x_matrix[155]) );
  DFFRHQX1 x_matrix_reg_2__7__10_ ( .D(n3809), .CK(clk), .RN(rst_n), .Q(
        x_matrix[458]) );
  DFFRHQX1 x_matrix_reg_6__3__10_ ( .D(n4257), .CK(clk), .RN(rst_n), .Q(
        x_matrix[154]) );
  DFFRHQX1 x_matrix_reg_2__7__0_ ( .D(n3819), .CK(clk), .RN(rst_n), .Q(
        x_matrix[448]) );
  DFFRHQX1 x_matrix_reg_6__3__0_ ( .D(n4267), .CK(clk), .RN(rst_n), .Q(
        x_matrix[144]) );
  DFFRHQX1 x_matrix_reg_3__7__9_ ( .D(n3938), .CK(clk), .RN(rst_n), .Q(
        x_matrix[361]) );
  DFFRHQX1 x_matrix_reg_7__3__9_ ( .D(n4386), .CK(clk), .RN(rst_n), .Q(
        x_matrix[73]) );
  DFFRHQX1 x_matrix_reg_3__7__8_ ( .D(n3939), .CK(clk), .RN(rst_n), .Q(
        x_matrix[360]) );
  DFFRHQX1 x_matrix_reg_7__3__8_ ( .D(n4387), .CK(clk), .RN(rst_n), .Q(
        x_matrix[72]) );
  DFFRHQX1 x_matrix_reg_3__7__7_ ( .D(n3940), .CK(clk), .RN(rst_n), .Q(
        x_matrix[359]) );
  DFFRHQX1 x_matrix_reg_7__3__7_ ( .D(n4388), .CK(clk), .RN(rst_n), .Q(
        x_matrix[71]) );
  DFFRHQX1 x_matrix_reg_3__7__6_ ( .D(n3941), .CK(clk), .RN(rst_n), .Q(
        x_matrix[358]) );
  DFFRHQX1 x_matrix_reg_7__3__6_ ( .D(n4389), .CK(clk), .RN(rst_n), .Q(
        x_matrix[70]) );
  DFFRHQX1 x_matrix_reg_5__0__15_ ( .D(n4076), .CK(clk), .RN(rst_n), .Q(
        x_matrix[255]) );
  DFFRHQX1 x_matrix_reg_7__4__15_ ( .D(n4396), .CK(clk), .RN(rst_n), .Q(
        x_matrix[63]) );
  DFFRHQX1 x_matrix_reg_5__0__14_ ( .D(n4077), .CK(clk), .RN(rst_n), .Q(
        x_matrix[254]) );
  DFFRHQX1 x_matrix_reg_7__4__14_ ( .D(n4397), .CK(clk), .RN(rst_n), .Q(
        x_matrix[62]) );
  DFFRHQX1 x_matrix_reg_5__0__13_ ( .D(n4078), .CK(clk), .RN(rst_n), .Q(
        x_matrix[253]) );
  DFFRHQX1 x_matrix_reg_7__4__13_ ( .D(n4398), .CK(clk), .RN(rst_n), .Q(
        x_matrix[61]) );
  DFFRHQX1 x_matrix_reg_5__0__12_ ( .D(n4079), .CK(clk), .RN(rst_n), .Q(
        x_matrix[252]) );
  DFFRHQX1 x_matrix_reg_7__4__12_ ( .D(n4399), .CK(clk), .RN(rst_n), .Q(
        x_matrix[60]) );
  DFFRHQX1 x_matrix_reg_3__7__5_ ( .D(n3942), .CK(clk), .RN(rst_n), .Q(
        x_matrix[357]) );
  DFFRHQX1 x_matrix_reg_7__3__5_ ( .D(n4390), .CK(clk), .RN(rst_n), .Q(
        x_matrix[69]) );
  DFFRHQX1 x_matrix_reg_5__0__11_ ( .D(n4080), .CK(clk), .RN(rst_n), .Q(
        x_matrix[251]) );
  DFFRHQX1 x_matrix_reg_7__4__11_ ( .D(n4400), .CK(clk), .RN(rst_n), .Q(
        x_matrix[59]) );
  DFFRHQX1 x_matrix_reg_5__0__10_ ( .D(n4081), .CK(clk), .RN(rst_n), .Q(
        x_matrix[250]) );
  DFFRHQX1 x_matrix_reg_7__4__10_ ( .D(n4401), .CK(clk), .RN(rst_n), .Q(
        x_matrix[58]) );
  DFFRHQX1 x_matrix_reg_5__0__9_ ( .D(n4082), .CK(clk), .RN(rst_n), .Q(
        x_matrix[249]) );
  DFFRHQX1 x_matrix_reg_7__4__9_ ( .D(n4402), .CK(clk), .RN(rst_n), .Q(
        x_matrix[57]) );
  DFFRHQX1 x_matrix_reg_5__0__8_ ( .D(n4083), .CK(clk), .RN(rst_n), .Q(
        x_matrix[248]) );
  DFFRHQX1 x_matrix_reg_7__4__8_ ( .D(n4403), .CK(clk), .RN(rst_n), .Q(
        x_matrix[56]) );
  DFFRHQX1 x_matrix_reg_5__0__7_ ( .D(n4084), .CK(clk), .RN(rst_n), .Q(
        x_matrix[247]) );
  DFFRHQX1 x_matrix_reg_7__4__7_ ( .D(n4404), .CK(clk), .RN(rst_n), .Q(
        x_matrix[55]) );
  DFFRHQX1 x_matrix_reg_5__0__6_ ( .D(n4085), .CK(clk), .RN(rst_n), .Q(
        x_matrix[246]) );
  DFFRHQX1 x_matrix_reg_7__4__6_ ( .D(n4405), .CK(clk), .RN(rst_n), .Q(
        x_matrix[54]) );
  DFFRHQX1 x_matrix_reg_5__0__5_ ( .D(n4086), .CK(clk), .RN(rst_n), .Q(
        x_matrix[245]) );
  DFFRHQX1 x_matrix_reg_7__4__5_ ( .D(n4406), .CK(clk), .RN(rst_n), .Q(
        x_matrix[53]) );
  DFFRHQX1 x_matrix_reg_5__0__4_ ( .D(n4087), .CK(clk), .RN(rst_n), .Q(
        x_matrix[244]) );
  DFFRHQX1 x_matrix_reg_7__4__4_ ( .D(n4407), .CK(clk), .RN(rst_n), .Q(
        x_matrix[52]) );
  DFFRHQX1 x_matrix_reg_5__0__3_ ( .D(n4088), .CK(clk), .RN(rst_n), .Q(
        x_matrix[243]) );
  DFFRHQX1 x_matrix_reg_7__4__3_ ( .D(n4408), .CK(clk), .RN(rst_n), .Q(
        x_matrix[51]) );
  DFFRHQX1 x_matrix_reg_5__0__2_ ( .D(n4089), .CK(clk), .RN(rst_n), .Q(
        x_matrix[242]) );
  DFFRHQX1 x_matrix_reg_7__4__2_ ( .D(n4409), .CK(clk), .RN(rst_n), .Q(
        x_matrix[50]) );
  DFFRHQX1 x_matrix_reg_3__7__4_ ( .D(n3943), .CK(clk), .RN(rst_n), .Q(
        x_matrix[356]) );
  DFFRHQX1 x_matrix_reg_7__3__4_ ( .D(n4391), .CK(clk), .RN(rst_n), .Q(
        x_matrix[68]) );
  DFFRHQX1 x_matrix_reg_5__0__1_ ( .D(n4090), .CK(clk), .RN(rst_n), .Q(
        x_matrix[241]) );
  DFFRHQX1 x_matrix_reg_7__4__1_ ( .D(n4410), .CK(clk), .RN(rst_n), .Q(
        x_matrix[49]) );
  DFFRHQX1 x_matrix_reg_5__0__0_ ( .D(n4091), .CK(clk), .RN(rst_n), .Q(
        x_matrix[240]) );
  DFFRHQX1 x_matrix_reg_7__4__0_ ( .D(n4411), .CK(clk), .RN(rst_n), .Q(
        x_matrix[48]) );
  DFFRHQX1 x_matrix_reg_1__5__15_ ( .D(n3644), .CK(clk), .RN(rst_n), .Q(
        x_matrix[575]) );
  DFFRHQX1 x_matrix_reg_5__1__15_ ( .D(n4092), .CK(clk), .RN(rst_n), .Q(
        x_matrix[239]) );
  DFFRHQX1 x_matrix_reg_1__5__14_ ( .D(n3645), .CK(clk), .RN(rst_n), .Q(
        x_matrix[574]) );
  DFFRHQX1 x_matrix_reg_5__1__14_ ( .D(n4093), .CK(clk), .RN(rst_n), .Q(
        x_matrix[238]) );
  DFFRHQX1 x_matrix_reg_1__5__13_ ( .D(n3646), .CK(clk), .RN(rst_n), .Q(
        x_matrix[573]) );
  DFFRHQX1 x_matrix_reg_5__1__13_ ( .D(n4094), .CK(clk), .RN(rst_n), .Q(
        x_matrix[237]) );
  DFFRHQX1 x_matrix_reg_1__5__12_ ( .D(n3647), .CK(clk), .RN(rst_n), .Q(
        x_matrix[572]) );
  DFFRHQX1 x_matrix_reg_5__1__12_ ( .D(n4095), .CK(clk), .RN(rst_n), .Q(
        x_matrix[236]) );
  DFFRHQX1 x_matrix_reg_1__5__11_ ( .D(n3648), .CK(clk), .RN(rst_n), .Q(
        x_matrix[571]) );
  DFFRHQX1 x_matrix_reg_5__1__11_ ( .D(n4096), .CK(clk), .RN(rst_n), .Q(
        x_matrix[235]) );
  DFFRHQX1 x_matrix_reg_1__5__10_ ( .D(n3649), .CK(clk), .RN(rst_n), .Q(
        x_matrix[570]) );
  DFFRHQX1 x_matrix_reg_5__1__10_ ( .D(n4097), .CK(clk), .RN(rst_n), .Q(
        x_matrix[234]) );
  DFFRHQX1 x_matrix_reg_1__5__9_ ( .D(n3650), .CK(clk), .RN(rst_n), .Q(
        x_matrix[569]) );
  DFFRHQX1 x_matrix_reg_5__1__9_ ( .D(n4098), .CK(clk), .RN(rst_n), .Q(
        x_matrix[233]) );
  DFFRHQX1 x_matrix_reg_1__5__8_ ( .D(n3651), .CK(clk), .RN(rst_n), .Q(
        x_matrix[568]) );
  DFFRHQX1 x_matrix_reg_5__1__8_ ( .D(n4099), .CK(clk), .RN(rst_n), .Q(
        x_matrix[232]) );
  DFFRHQX1 x_matrix_reg_3__7__3_ ( .D(n3944), .CK(clk), .RN(rst_n), .Q(
        x_matrix[355]) );
  DFFRHQX1 x_matrix_reg_7__3__3_ ( .D(n4392), .CK(clk), .RN(rst_n), .Q(
        x_matrix[67]) );
  DFFRHQX1 x_matrix_reg_1__5__7_ ( .D(n3652), .CK(clk), .RN(rst_n), .Q(
        x_matrix[567]) );
  DFFRHQX1 x_matrix_reg_5__1__7_ ( .D(n4100), .CK(clk), .RN(rst_n), .Q(
        x_matrix[231]) );
  DFFRHQX1 x_matrix_reg_1__5__6_ ( .D(n3653), .CK(clk), .RN(rst_n), .Q(
        x_matrix[566]) );
  DFFRHQX1 x_matrix_reg_5__1__6_ ( .D(n4101), .CK(clk), .RN(rst_n), .Q(
        x_matrix[230]) );
  DFFRHQX1 x_matrix_reg_1__5__5_ ( .D(n3654), .CK(clk), .RN(rst_n), .Q(
        x_matrix[565]) );
  DFFRHQX1 x_matrix_reg_5__1__5_ ( .D(n4102), .CK(clk), .RN(rst_n), .Q(
        x_matrix[229]) );
  DFFRHQX1 x_matrix_reg_1__5__4_ ( .D(n3655), .CK(clk), .RN(rst_n), .Q(
        x_matrix[564]) );
  DFFRHQX1 x_matrix_reg_5__1__4_ ( .D(n4103), .CK(clk), .RN(rst_n), .Q(
        x_matrix[228]) );
  DFFRHQX1 x_matrix_reg_1__5__3_ ( .D(n3656), .CK(clk), .RN(rst_n), .Q(
        x_matrix[563]) );
  DFFRHQX1 x_matrix_reg_5__1__3_ ( .D(n4104), .CK(clk), .RN(rst_n), .Q(
        x_matrix[227]) );
  DFFRHQX1 x_matrix_reg_1__5__2_ ( .D(n3657), .CK(clk), .RN(rst_n), .Q(
        x_matrix[562]) );
  DFFRHQX1 x_matrix_reg_5__1__2_ ( .D(n4105), .CK(clk), .RN(rst_n), .Q(
        x_matrix[226]) );
  DFFRHQX1 x_matrix_reg_1__5__1_ ( .D(n3658), .CK(clk), .RN(rst_n), .Q(
        x_matrix[561]) );
  DFFRHQX1 x_matrix_reg_5__1__1_ ( .D(n4106), .CK(clk), .RN(rst_n), .Q(
        x_matrix[225]) );
  DFFRHQX1 x_matrix_reg_1__5__0_ ( .D(n3659), .CK(clk), .RN(rst_n), .Q(
        x_matrix[560]) );
  DFFRHQX1 x_matrix_reg_5__1__0_ ( .D(n4107), .CK(clk), .RN(rst_n), .Q(
        x_matrix[224]) );
  DFFRHQX1 x_matrix_reg_1__6__15_ ( .D(n3660), .CK(clk), .RN(rst_n), .Q(
        x_matrix[559]) );
  DFFRHQX1 x_matrix_reg_5__2__15_ ( .D(n4108), .CK(clk), .RN(rst_n), .Q(
        x_matrix[223]) );
  DFFRHQX1 x_matrix_reg_1__6__14_ ( .D(n3661), .CK(clk), .RN(rst_n), .Q(
        x_matrix[558]) );
  DFFRHQX1 x_matrix_reg_5__2__14_ ( .D(n4109), .CK(clk), .RN(rst_n), .Q(
        x_matrix[222]) );
  DFFRHQX1 x_matrix_reg_3__7__2_ ( .D(n3945), .CK(clk), .RN(rst_n), .Q(
        x_matrix[354]) );
  DFFRHQX1 x_matrix_reg_7__3__2_ ( .D(n4393), .CK(clk), .RN(rst_n), .Q(
        x_matrix[66]) );
  DFFRHQX1 x_matrix_reg_1__6__13_ ( .D(n3662), .CK(clk), .RN(rst_n), .Q(
        x_matrix[557]) );
  DFFRHQX1 x_matrix_reg_5__2__13_ ( .D(n4110), .CK(clk), .RN(rst_n), .Q(
        x_matrix[221]) );
  DFFRHQX1 x_matrix_reg_1__6__12_ ( .D(n3663), .CK(clk), .RN(rst_n), .Q(
        x_matrix[556]) );
  DFFRHQX1 x_matrix_reg_5__2__12_ ( .D(n4111), .CK(clk), .RN(rst_n), .Q(
        x_matrix[220]) );
  DFFRHQX1 x_matrix_reg_1__6__11_ ( .D(n3664), .CK(clk), .RN(rst_n), .Q(
        x_matrix[555]) );
  DFFRHQX1 x_matrix_reg_5__2__11_ ( .D(n4112), .CK(clk), .RN(rst_n), .Q(
        x_matrix[219]) );
  DFFRHQX1 x_matrix_reg_1__6__10_ ( .D(n3665), .CK(clk), .RN(rst_n), .Q(
        x_matrix[554]) );
  DFFRHQX1 x_matrix_reg_5__2__10_ ( .D(n4113), .CK(clk), .RN(rst_n), .Q(
        x_matrix[218]) );
  DFFRHQX1 x_matrix_reg_1__6__9_ ( .D(n3666), .CK(clk), .RN(rst_n), .Q(
        x_matrix[553]) );
  DFFRHQX1 x_matrix_reg_5__2__9_ ( .D(n4114), .CK(clk), .RN(rst_n), .Q(
        x_matrix[217]) );
  DFFRHQX1 x_matrix_reg_1__6__8_ ( .D(n3667), .CK(clk), .RN(rst_n), .Q(
        x_matrix[552]) );
  DFFRHQX1 x_matrix_reg_5__2__8_ ( .D(n4115), .CK(clk), .RN(rst_n), .Q(
        x_matrix[216]) );
  DFFRHQX1 x_matrix_reg_1__6__7_ ( .D(n3668), .CK(clk), .RN(rst_n), .Q(
        x_matrix[551]) );
  DFFRHQX1 x_matrix_reg_5__2__7_ ( .D(n4116), .CK(clk), .RN(rst_n), .Q(
        x_matrix[215]) );
  DFFRHQX1 x_matrix_reg_1__6__6_ ( .D(n3669), .CK(clk), .RN(rst_n), .Q(
        x_matrix[550]) );
  DFFRHQX1 x_matrix_reg_5__2__6_ ( .D(n4117), .CK(clk), .RN(rst_n), .Q(
        x_matrix[214]) );
  DFFRHQX1 x_matrix_reg_1__6__5_ ( .D(n3670), .CK(clk), .RN(rst_n), .Q(
        x_matrix[549]) );
  DFFRHQX1 x_matrix_reg_5__2__5_ ( .D(n4118), .CK(clk), .RN(rst_n), .Q(
        x_matrix[213]) );
  DFFRHQX1 x_matrix_reg_1__6__4_ ( .D(n3671), .CK(clk), .RN(rst_n), .Q(
        x_matrix[548]) );
  DFFRHQX1 x_matrix_reg_5__2__4_ ( .D(n4119), .CK(clk), .RN(rst_n), .Q(
        x_matrix[212]) );
  DFFRHQX1 x_matrix_reg_3__7__1_ ( .D(n3946), .CK(clk), .RN(rst_n), .Q(
        x_matrix[353]) );
  DFFRHQX1 x_matrix_reg_7__3__1_ ( .D(n4394), .CK(clk), .RN(rst_n), .Q(
        x_matrix[65]) );
  DFFRHQX1 x_matrix_reg_1__6__3_ ( .D(n3672), .CK(clk), .RN(rst_n), .Q(
        x_matrix[547]) );
  DFFRHQX1 x_matrix_reg_5__2__3_ ( .D(n4120), .CK(clk), .RN(rst_n), .Q(
        x_matrix[211]) );
  DFFRHQX1 x_matrix_reg_1__6__2_ ( .D(n3673), .CK(clk), .RN(rst_n), .Q(
        x_matrix[546]) );
  DFFRHQX1 x_matrix_reg_5__2__2_ ( .D(n4121), .CK(clk), .RN(rst_n), .Q(
        x_matrix[210]) );
  DFFRHQX1 x_matrix_reg_1__6__1_ ( .D(n3674), .CK(clk), .RN(rst_n), .Q(
        x_matrix[545]) );
  DFFRHQX1 x_matrix_reg_5__2__1_ ( .D(n4122), .CK(clk), .RN(rst_n), .Q(
        x_matrix[209]) );
  DFFRHQX1 x_matrix_reg_1__6__0_ ( .D(n3675), .CK(clk), .RN(rst_n), .Q(
        x_matrix[544]) );
  DFFRHQX1 x_matrix_reg_5__2__0_ ( .D(n4123), .CK(clk), .RN(rst_n), .Q(
        x_matrix[208]) );
  DFFRHQX1 x_matrix_reg_3__7__15_ ( .D(n3932), .CK(clk), .RN(rst_n), .Q(
        x_matrix[367]) );
  DFFRHQX1 x_matrix_reg_7__3__15_ ( .D(n4380), .CK(clk), .RN(rst_n), .Q(
        x_matrix[79]) );
  DFFRHQX1 x_matrix_reg_3__7__14_ ( .D(n3933), .CK(clk), .RN(rst_n), .Q(
        x_matrix[366]) );
  DFFRHQX1 x_matrix_reg_7__3__14_ ( .D(n4381), .CK(clk), .RN(rst_n), .Q(
        x_matrix[78]) );
  DFFRHQX1 x_matrix_reg_3__7__13_ ( .D(n3934), .CK(clk), .RN(rst_n), .Q(
        x_matrix[365]) );
  DFFRHQX1 x_matrix_reg_7__3__13_ ( .D(n4382), .CK(clk), .RN(rst_n), .Q(
        x_matrix[77]) );
  DFFRHQX1 x_matrix_reg_3__7__12_ ( .D(n3935), .CK(clk), .RN(rst_n), .Q(
        x_matrix[364]) );
  DFFRHQX1 x_matrix_reg_7__3__12_ ( .D(n4383), .CK(clk), .RN(rst_n), .Q(
        x_matrix[76]) );
  DFFRHQX1 x_matrix_reg_3__7__11_ ( .D(n3936), .CK(clk), .RN(rst_n), .Q(
        x_matrix[363]) );
  DFFRHQX1 x_matrix_reg_7__3__11_ ( .D(n4384), .CK(clk), .RN(rst_n), .Q(
        x_matrix[75]) );
  DFFRHQX1 x_matrix_reg_3__7__10_ ( .D(n3937), .CK(clk), .RN(rst_n), .Q(
        x_matrix[362]) );
  DFFRHQX1 x_matrix_reg_7__3__10_ ( .D(n4385), .CK(clk), .RN(rst_n), .Q(
        x_matrix[74]) );
  DFFRHQX1 x_matrix_reg_3__7__0_ ( .D(n3947), .CK(clk), .RN(rst_n), .Q(
        x_matrix[352]) );
  DFFRHQX1 x_matrix_reg_7__3__0_ ( .D(n4395), .CK(clk), .RN(rst_n), .Q(
        x_matrix[64]) );
  DFFRHQX1 cal_out_reg_5__32_ ( .D(n2019), .CK(clk), .RN(rst_n), .Q(
        cal_out[392]) );
  DFFRHQX1 cal_out_reg_11__32_ ( .D(n2259), .CK(clk), .RN(rst_n), .Q(
        cal_out[152]) );
  DFFRHQX1 cal_out_reg_4__32_ ( .D(n1979), .CK(clk), .RN(rst_n), .Q(
        cal_out[432]) );
  DFFRHQX1 cal_out_reg_6__32_ ( .D(n2059), .CK(clk), .RN(rst_n), .Q(
        cal_out[352]) );
  DFFRHQX1 length_reg_reg_4__5_ ( .D(n1746), .CK(clk), .RN(rst_n), .Q(
        length_reg[65]) );
  DFFRHQX1 length_reg_reg_6__5_ ( .D(n1758), .CK(clk), .RN(rst_n), .Q(
        length_reg[53]) );
  DFFRHQX1 cal_out_reg_10__32_ ( .D(n2219), .CK(clk), .RN(rst_n), .Q(
        cal_out[192]) );
  DFFRX1 x_matrix_reg_1__7__9_ ( .D(n3682), .CK(clk), .RN(rst_n), .QN(n424) );
  DFFRX1 x_matrix_reg_5__3__9_ ( .D(n4130), .CK(clk), .RN(rst_n), .QN(n536) );
  DFFRX1 x_matrix_reg_1__7__8_ ( .D(n3683), .CK(clk), .RN(rst_n), .QN(n425) );
  DFFRX1 x_matrix_reg_5__3__8_ ( .D(n4131), .CK(clk), .RN(rst_n), .QN(n537) );
  DFFRX1 x_matrix_reg_1__7__7_ ( .D(n3684), .CK(clk), .RN(rst_n), .QN(n426) );
  DFFRX1 x_matrix_reg_5__3__7_ ( .D(n4132), .CK(clk), .RN(rst_n), .QN(n538) );
  DFFRX1 x_matrix_reg_1__7__6_ ( .D(n3685), .CK(clk), .RN(rst_n), .QN(n427) );
  DFFRX1 x_matrix_reg_5__3__6_ ( .D(n4133), .CK(clk), .RN(rst_n), .QN(n539) );
  DFFRX1 x_matrix_reg_5__4__15_ ( .D(n4140), .CK(clk), .RN(rst_n), .QN(n546)
         );
  DFFRX1 x_matrix_reg_7__0__15_ ( .D(n4332), .CK(clk), .RN(rst_n), .QN(n610)
         );
  DFFRX1 x_matrix_reg_5__4__14_ ( .D(n4141), .CK(clk), .RN(rst_n), .QN(n547)
         );
  DFFRX1 x_matrix_reg_7__0__14_ ( .D(n4333), .CK(clk), .RN(rst_n), .QN(n611)
         );
  DFFRX1 x_matrix_reg_5__4__13_ ( .D(n4142), .CK(clk), .RN(rst_n), .QN(n548)
         );
  DFFRX1 x_matrix_reg_7__0__13_ ( .D(n4334), .CK(clk), .RN(rst_n), .QN(n612)
         );
  DFFRX1 x_matrix_reg_5__4__12_ ( .D(n4143), .CK(clk), .RN(rst_n), .QN(n549)
         );
  DFFRX1 x_matrix_reg_7__0__12_ ( .D(n4335), .CK(clk), .RN(rst_n), .QN(n613)
         );
  DFFRX1 x_matrix_reg_1__7__5_ ( .D(n3686), .CK(clk), .RN(rst_n), .QN(n428) );
  DFFRX1 x_matrix_reg_5__3__5_ ( .D(n4134), .CK(clk), .RN(rst_n), .QN(n540) );
  DFFRX1 x_matrix_reg_5__4__11_ ( .D(n4144), .CK(clk), .RN(rst_n), .QN(n550)
         );
  DFFRX1 x_matrix_reg_7__0__11_ ( .D(n4336), .CK(clk), .RN(rst_n), .QN(n614)
         );
  DFFRX1 x_matrix_reg_5__4__10_ ( .D(n4145), .CK(clk), .RN(rst_n), .QN(n551)
         );
  DFFRX1 x_matrix_reg_7__0__10_ ( .D(n4337), .CK(clk), .RN(rst_n), .QN(n615)
         );
  DFFRX1 x_matrix_reg_5__4__9_ ( .D(n4146), .CK(clk), .RN(rst_n), .QN(n552) );
  DFFRX1 x_matrix_reg_7__0__9_ ( .D(n4338), .CK(clk), .RN(rst_n), .QN(n616) );
  DFFRX1 x_matrix_reg_5__4__8_ ( .D(n4147), .CK(clk), .RN(rst_n), .QN(n553) );
  DFFRX1 x_matrix_reg_7__0__8_ ( .D(n4339), .CK(clk), .RN(rst_n), .QN(n617) );
  DFFRX1 x_matrix_reg_5__4__7_ ( .D(n4148), .CK(clk), .RN(rst_n), .QN(n554) );
  DFFRX1 x_matrix_reg_7__0__7_ ( .D(n4340), .CK(clk), .RN(rst_n), .QN(n618) );
  DFFRX1 x_matrix_reg_5__4__6_ ( .D(n4149), .CK(clk), .RN(rst_n), .QN(n555) );
  DFFRX1 x_matrix_reg_7__0__6_ ( .D(n4341), .CK(clk), .RN(rst_n), .QN(n619) );
  DFFRX1 x_matrix_reg_5__4__5_ ( .D(n4150), .CK(clk), .RN(rst_n), .QN(n556) );
  DFFRX1 x_matrix_reg_7__0__5_ ( .D(n4342), .CK(clk), .RN(rst_n), .QN(n620) );
  DFFRX1 x_matrix_reg_5__4__4_ ( .D(n4151), .CK(clk), .RN(rst_n), .QN(n557) );
  DFFRX1 x_matrix_reg_7__0__4_ ( .D(n4343), .CK(clk), .RN(rst_n), .QN(n621) );
  DFFRX1 x_matrix_reg_5__4__3_ ( .D(n4152), .CK(clk), .RN(rst_n), .QN(n558) );
  DFFRX1 x_matrix_reg_7__0__3_ ( .D(n4344), .CK(clk), .RN(rst_n), .QN(n622) );
  DFFRX1 x_matrix_reg_5__4__2_ ( .D(n4153), .CK(clk), .RN(rst_n), .QN(n559) );
  DFFRX1 x_matrix_reg_7__0__2_ ( .D(n4345), .CK(clk), .RN(rst_n), .QN(n623) );
  DFFRX1 x_matrix_reg_1__7__4_ ( .D(n3687), .CK(clk), .RN(rst_n), .QN(n429) );
  DFFRX1 x_matrix_reg_5__3__4_ ( .D(n4135), .CK(clk), .RN(rst_n), .QN(n541) );
  DFFRX1 x_matrix_reg_5__4__1_ ( .D(n4154), .CK(clk), .RN(rst_n), .QN(n560) );
  DFFRX1 x_matrix_reg_7__0__1_ ( .D(n4346), .CK(clk), .RN(rst_n), .QN(n624) );
  DFFRX1 x_matrix_reg_5__4__0_ ( .D(n4155), .CK(clk), .RN(rst_n), .QN(n561) );
  DFFRX1 x_matrix_reg_7__0__0_ ( .D(n4347), .CK(clk), .RN(rst_n), .QN(n625) );
  DFFRX1 x_matrix_reg_3__5__15_ ( .D(n3900), .CK(clk), .RN(rst_n), .QN(n466)
         );
  DFFRX1 x_matrix_reg_7__1__15_ ( .D(n4348), .CK(clk), .RN(rst_n), .QN(n626)
         );
  DFFRX1 x_matrix_reg_3__5__14_ ( .D(n3901), .CK(clk), .RN(rst_n), .QN(n467)
         );
  DFFRX1 x_matrix_reg_7__1__14_ ( .D(n4349), .CK(clk), .RN(rst_n), .QN(n627)
         );
  DFFRX1 x_matrix_reg_3__5__13_ ( .D(n3902), .CK(clk), .RN(rst_n), .QN(n468)
         );
  DFFRX1 x_matrix_reg_7__1__13_ ( .D(n4350), .CK(clk), .RN(rst_n), .QN(n628)
         );
  DFFRX1 x_matrix_reg_3__5__12_ ( .D(n3903), .CK(clk), .RN(rst_n), .QN(n469)
         );
  DFFRX1 x_matrix_reg_7__1__12_ ( .D(n4351), .CK(clk), .RN(rst_n), .QN(n629)
         );
  DFFRX1 x_matrix_reg_3__5__11_ ( .D(n3904), .CK(clk), .RN(rst_n), .QN(n470)
         );
  DFFRX1 x_matrix_reg_7__1__11_ ( .D(n4352), .CK(clk), .RN(rst_n), .QN(n630)
         );
  DFFRX1 x_matrix_reg_3__5__10_ ( .D(n3905), .CK(clk), .RN(rst_n), .QN(n471)
         );
  DFFRX1 x_matrix_reg_7__1__10_ ( .D(n4353), .CK(clk), .RN(rst_n), .QN(n631)
         );
  DFFRX1 x_matrix_reg_3__5__9_ ( .D(n3906), .CK(clk), .RN(rst_n), .QN(n472) );
  DFFRX1 x_matrix_reg_7__1__9_ ( .D(n4354), .CK(clk), .RN(rst_n), .QN(n632) );
  DFFRX1 x_matrix_reg_3__5__8_ ( .D(n3907), .CK(clk), .RN(rst_n), .QN(n473) );
  DFFRX1 x_matrix_reg_7__1__8_ ( .D(n4355), .CK(clk), .RN(rst_n), .QN(n633) );
  DFFRX1 x_matrix_reg_1__7__3_ ( .D(n3688), .CK(clk), .RN(rst_n), .QN(n430) );
  DFFRX1 x_matrix_reg_5__3__3_ ( .D(n4136), .CK(clk), .RN(rst_n), .QN(n542) );
  DFFRX1 x_matrix_reg_3__5__7_ ( .D(n3908), .CK(clk), .RN(rst_n), .QN(n474) );
  DFFRX1 x_matrix_reg_7__1__7_ ( .D(n4356), .CK(clk), .RN(rst_n), .QN(n634) );
  DFFRX1 x_matrix_reg_3__5__6_ ( .D(n3909), .CK(clk), .RN(rst_n), .QN(n475) );
  DFFRX1 x_matrix_reg_7__1__6_ ( .D(n4357), .CK(clk), .RN(rst_n), .QN(n635) );
  DFFRX1 x_matrix_reg_3__5__5_ ( .D(n3910), .CK(clk), .RN(rst_n), .QN(n476) );
  DFFRX1 x_matrix_reg_7__1__5_ ( .D(n4358), .CK(clk), .RN(rst_n), .QN(n636) );
  DFFRX1 x_matrix_reg_3__5__4_ ( .D(n3911), .CK(clk), .RN(rst_n), .QN(n477) );
  DFFRX1 x_matrix_reg_7__1__4_ ( .D(n4359), .CK(clk), .RN(rst_n), .QN(n637) );
  DFFRX1 x_matrix_reg_3__5__3_ ( .D(n3912), .CK(clk), .RN(rst_n), .QN(n478) );
  DFFRX1 x_matrix_reg_7__1__3_ ( .D(n4360), .CK(clk), .RN(rst_n), .QN(n638) );
  DFFRX1 x_matrix_reg_3__5__2_ ( .D(n3913), .CK(clk), .RN(rst_n), .QN(n479) );
  DFFRX1 x_matrix_reg_7__1__2_ ( .D(n4361), .CK(clk), .RN(rst_n), .QN(n639) );
  DFFRX1 x_matrix_reg_3__5__1_ ( .D(n3914), .CK(clk), .RN(rst_n), .QN(n480) );
  DFFRX1 x_matrix_reg_7__1__1_ ( .D(n4362), .CK(clk), .RN(rst_n), .QN(n640) );
  DFFRX1 x_matrix_reg_3__5__0_ ( .D(n3915), .CK(clk), .RN(rst_n), .QN(n481) );
  DFFRX1 x_matrix_reg_7__1__0_ ( .D(n4363), .CK(clk), .RN(rst_n), .QN(n641) );
  DFFRX1 x_matrix_reg_3__6__15_ ( .D(n3916), .CK(clk), .RN(rst_n), .QN(n482)
         );
  DFFRX1 x_matrix_reg_7__2__15_ ( .D(n4364), .CK(clk), .RN(rst_n), .QN(n642)
         );
  DFFRX1 x_matrix_reg_3__6__14_ ( .D(n3917), .CK(clk), .RN(rst_n), .QN(n483)
         );
  DFFRX1 x_matrix_reg_7__2__14_ ( .D(n4365), .CK(clk), .RN(rst_n), .QN(n643)
         );
  DFFRX1 x_matrix_reg_1__7__2_ ( .D(n3689), .CK(clk), .RN(rst_n), .QN(n431) );
  DFFRX1 x_matrix_reg_5__3__2_ ( .D(n4137), .CK(clk), .RN(rst_n), .QN(n543) );
  DFFRX1 x_matrix_reg_3__6__13_ ( .D(n3918), .CK(clk), .RN(rst_n), .QN(n484)
         );
  DFFRX1 x_matrix_reg_7__2__13_ ( .D(n4366), .CK(clk), .RN(rst_n), .QN(n644)
         );
  DFFRX1 x_matrix_reg_3__6__12_ ( .D(n3919), .CK(clk), .RN(rst_n), .QN(n485)
         );
  DFFRX1 x_matrix_reg_7__2__12_ ( .D(n4367), .CK(clk), .RN(rst_n), .QN(n645)
         );
  DFFRX1 x_matrix_reg_3__6__11_ ( .D(n3920), .CK(clk), .RN(rst_n), .QN(n486)
         );
  DFFRX1 x_matrix_reg_7__2__11_ ( .D(n4368), .CK(clk), .RN(rst_n), .QN(n646)
         );
  DFFRX1 x_matrix_reg_3__6__10_ ( .D(n3921), .CK(clk), .RN(rst_n), .QN(n487)
         );
  DFFRX1 x_matrix_reg_7__2__10_ ( .D(n4369), .CK(clk), .RN(rst_n), .QN(n647)
         );
  DFFRX1 x_matrix_reg_3__6__9_ ( .D(n3922), .CK(clk), .RN(rst_n), .QN(n488) );
  DFFRX1 x_matrix_reg_7__2__9_ ( .D(n4370), .CK(clk), .RN(rst_n), .QN(n648) );
  DFFRX1 x_matrix_reg_3__6__8_ ( .D(n3923), .CK(clk), .RN(rst_n), .QN(n489) );
  DFFRX1 x_matrix_reg_7__2__8_ ( .D(n4371), .CK(clk), .RN(rst_n), .QN(n649) );
  DFFRX1 x_matrix_reg_3__6__7_ ( .D(n3924), .CK(clk), .RN(rst_n), .QN(n490) );
  DFFRX1 x_matrix_reg_7__2__7_ ( .D(n4372), .CK(clk), .RN(rst_n), .QN(n650) );
  DFFRX1 x_matrix_reg_3__6__6_ ( .D(n3925), .CK(clk), .RN(rst_n), .QN(n491) );
  DFFRX1 x_matrix_reg_7__2__6_ ( .D(n4373), .CK(clk), .RN(rst_n), .QN(n651) );
  DFFRX1 x_matrix_reg_3__6__5_ ( .D(n3926), .CK(clk), .RN(rst_n), .QN(n492) );
  DFFRX1 x_matrix_reg_7__2__5_ ( .D(n4374), .CK(clk), .RN(rst_n), .QN(n652) );
  DFFRX1 x_matrix_reg_3__6__4_ ( .D(n3927), .CK(clk), .RN(rst_n), .QN(n493) );
  DFFRX1 x_matrix_reg_7__2__4_ ( .D(n4375), .CK(clk), .RN(rst_n), .QN(n653) );
  DFFRX1 x_matrix_reg_1__7__1_ ( .D(n3690), .CK(clk), .RN(rst_n), .QN(n432) );
  DFFRX1 x_matrix_reg_5__3__1_ ( .D(n4138), .CK(clk), .RN(rst_n), .QN(n544) );
  DFFRX1 x_matrix_reg_3__6__3_ ( .D(n3928), .CK(clk), .RN(rst_n), .QN(n494) );
  DFFRX1 x_matrix_reg_7__2__3_ ( .D(n4376), .CK(clk), .RN(rst_n), .QN(n654) );
  DFFRX1 x_matrix_reg_3__6__2_ ( .D(n3929), .CK(clk), .RN(rst_n), .QN(n495) );
  DFFRX1 x_matrix_reg_7__2__2_ ( .D(n4377), .CK(clk), .RN(rst_n), .QN(n655) );
  DFFRX1 x_matrix_reg_3__6__1_ ( .D(n3930), .CK(clk), .RN(rst_n), .QN(n496) );
  DFFRX1 x_matrix_reg_7__2__1_ ( .D(n4378), .CK(clk), .RN(rst_n), .QN(n656) );
  DFFRX1 x_matrix_reg_3__6__0_ ( .D(n3931), .CK(clk), .RN(rst_n), .QN(n497) );
  DFFRX1 x_matrix_reg_7__2__0_ ( .D(n4379), .CK(clk), .RN(rst_n), .QN(n657) );
  DFFRX1 x_matrix_reg_1__7__15_ ( .D(n3676), .CK(clk), .RN(rst_n), .QN(n418)
         );
  DFFRX1 x_matrix_reg_5__3__15_ ( .D(n4124), .CK(clk), .RN(rst_n), .QN(n530)
         );
  DFFRX1 x_matrix_reg_1__7__14_ ( .D(n3677), .CK(clk), .RN(rst_n), .QN(n419)
         );
  DFFRX1 x_matrix_reg_5__3__14_ ( .D(n4125), .CK(clk), .RN(rst_n), .QN(n531)
         );
  DFFRX1 x_matrix_reg_1__7__13_ ( .D(n3678), .CK(clk), .RN(rst_n), .QN(n420)
         );
  DFFRX1 x_matrix_reg_5__3__13_ ( .D(n4126), .CK(clk), .RN(rst_n), .QN(n532)
         );
  DFFRX1 x_matrix_reg_1__7__12_ ( .D(n3679), .CK(clk), .RN(rst_n), .QN(n421)
         );
  DFFRX1 x_matrix_reg_5__3__12_ ( .D(n4127), .CK(clk), .RN(rst_n), .QN(n533)
         );
  DFFRX1 x_matrix_reg_1__7__11_ ( .D(n3680), .CK(clk), .RN(rst_n), .QN(n422)
         );
  DFFRX1 x_matrix_reg_5__3__11_ ( .D(n4128), .CK(clk), .RN(rst_n), .QN(n534)
         );
  DFFRX1 x_matrix_reg_1__7__10_ ( .D(n3681), .CK(clk), .RN(rst_n), .QN(n423)
         );
  DFFRX1 x_matrix_reg_5__3__10_ ( .D(n4129), .CK(clk), .RN(rst_n), .QN(n535)
         );
  DFFRX1 x_matrix_reg_1__7__0_ ( .D(n3691), .CK(clk), .RN(rst_n), .QN(n433) );
  DFFRX1 x_matrix_reg_5__3__0_ ( .D(n4139), .CK(clk), .RN(rst_n), .QN(n545) );
  DFFRX1 x_matrix_reg_0__7__9_ ( .D(n3554), .CK(clk), .RN(rst_n), .QN(n376) );
  DFFRX1 x_matrix_reg_4__3__9_ ( .D(n4002), .CK(clk), .RN(rst_n), .QN(n504) );
  DFFRX1 x_matrix_reg_0__7__8_ ( .D(n3555), .CK(clk), .RN(rst_n), .QN(n377) );
  DFFRX1 x_matrix_reg_4__3__8_ ( .D(n4003), .CK(clk), .RN(rst_n), .QN(n505) );
  DFFRX1 x_matrix_reg_0__7__7_ ( .D(n3556), .CK(clk), .RN(rst_n), .QN(n378) );
  DFFRX1 x_matrix_reg_4__3__7_ ( .D(n4004), .CK(clk), .RN(rst_n), .QN(n506) );
  DFFRX1 x_matrix_reg_0__7__6_ ( .D(n3557), .CK(clk), .RN(rst_n), .QN(n379) );
  DFFRX1 x_matrix_reg_4__3__6_ ( .D(n4005), .CK(clk), .RN(rst_n), .QN(n507) );
  DFFRX1 x_matrix_reg_4__4__15_ ( .D(n4012), .CK(clk), .RN(rst_n), .QN(n514)
         );
  DFFRX1 x_matrix_reg_6__0__15_ ( .D(n4204), .CK(clk), .RN(rst_n), .QN(n562)
         );
  DFFRX1 x_matrix_reg_4__4__14_ ( .D(n4013), .CK(clk), .RN(rst_n), .QN(n515)
         );
  DFFRX1 x_matrix_reg_6__0__14_ ( .D(n4205), .CK(clk), .RN(rst_n), .QN(n563)
         );
  DFFRX1 x_matrix_reg_4__4__13_ ( .D(n4014), .CK(clk), .RN(rst_n), .QN(n516)
         );
  DFFRX1 x_matrix_reg_6__0__13_ ( .D(n4206), .CK(clk), .RN(rst_n), .QN(n564)
         );
  DFFRX1 x_matrix_reg_4__4__12_ ( .D(n4015), .CK(clk), .RN(rst_n), .QN(n517)
         );
  DFFRX1 x_matrix_reg_6__0__12_ ( .D(n4207), .CK(clk), .RN(rst_n), .QN(n565)
         );
  DFFRX1 x_matrix_reg_0__7__5_ ( .D(n3558), .CK(clk), .RN(rst_n), .QN(n380) );
  DFFRX1 x_matrix_reg_4__3__5_ ( .D(n4006), .CK(clk), .RN(rst_n), .QN(n508) );
  DFFRX1 x_matrix_reg_4__4__11_ ( .D(n4016), .CK(clk), .RN(rst_n), .QN(n518)
         );
  DFFRX1 x_matrix_reg_6__0__11_ ( .D(n4208), .CK(clk), .RN(rst_n), .QN(n566)
         );
  DFFRX1 x_matrix_reg_4__4__10_ ( .D(n4017), .CK(clk), .RN(rst_n), .QN(n519)
         );
  DFFRX1 x_matrix_reg_6__0__10_ ( .D(n4209), .CK(clk), .RN(rst_n), .QN(n567)
         );
  DFFRX1 x_matrix_reg_4__4__9_ ( .D(n4018), .CK(clk), .RN(rst_n), .QN(n520) );
  DFFRX1 x_matrix_reg_6__0__9_ ( .D(n4210), .CK(clk), .RN(rst_n), .QN(n568) );
  DFFRX1 x_matrix_reg_4__4__8_ ( .D(n4019), .CK(clk), .RN(rst_n), .QN(n521) );
  DFFRX1 x_matrix_reg_6__0__8_ ( .D(n4211), .CK(clk), .RN(rst_n), .QN(n569) );
  DFFRX1 x_matrix_reg_4__4__7_ ( .D(n4020), .CK(clk), .RN(rst_n), .QN(n522) );
  DFFRX1 x_matrix_reg_6__0__7_ ( .D(n4212), .CK(clk), .RN(rst_n), .QN(n570) );
  DFFRX1 x_matrix_reg_4__4__6_ ( .D(n4021), .CK(clk), .RN(rst_n), .QN(n523) );
  DFFRX1 x_matrix_reg_6__0__6_ ( .D(n4213), .CK(clk), .RN(rst_n), .QN(n571) );
  DFFRX1 x_matrix_reg_4__4__5_ ( .D(n4022), .CK(clk), .RN(rst_n), .QN(n524) );
  DFFRX1 x_matrix_reg_6__0__5_ ( .D(n4214), .CK(clk), .RN(rst_n), .QN(n572) );
  DFFRX1 x_matrix_reg_4__4__4_ ( .D(n4023), .CK(clk), .RN(rst_n), .QN(n525) );
  DFFRX1 x_matrix_reg_6__0__4_ ( .D(n4215), .CK(clk), .RN(rst_n), .QN(n573) );
  DFFRX1 x_matrix_reg_4__4__3_ ( .D(n4024), .CK(clk), .RN(rst_n), .QN(n526) );
  DFFRX1 x_matrix_reg_6__0__3_ ( .D(n4216), .CK(clk), .RN(rst_n), .QN(n574) );
  DFFRX1 x_matrix_reg_4__4__2_ ( .D(n4025), .CK(clk), .RN(rst_n), .QN(n527) );
  DFFRX1 x_matrix_reg_6__0__2_ ( .D(n4217), .CK(clk), .RN(rst_n), .QN(n575) );
  DFFRX1 x_matrix_reg_0__7__4_ ( .D(n3559), .CK(clk), .RN(rst_n), .QN(n381) );
  DFFRX1 x_matrix_reg_4__3__4_ ( .D(n4007), .CK(clk), .RN(rst_n), .QN(n509) );
  DFFRX1 x_matrix_reg_4__4__1_ ( .D(n4026), .CK(clk), .RN(rst_n), .QN(n528) );
  DFFRX1 x_matrix_reg_6__0__1_ ( .D(n4218), .CK(clk), .RN(rst_n), .QN(n576) );
  DFFRX1 x_matrix_reg_4__4__0_ ( .D(n4027), .CK(clk), .RN(rst_n), .QN(n529) );
  DFFRX1 x_matrix_reg_6__0__0_ ( .D(n4219), .CK(clk), .RN(rst_n), .QN(n577) );
  DFFRX1 x_matrix_reg_2__5__15_ ( .D(n3772), .CK(clk), .RN(rst_n), .QN(n434)
         );
  DFFRX1 x_matrix_reg_6__1__15_ ( .D(n4220), .CK(clk), .RN(rst_n), .QN(n578)
         );
  DFFRX1 x_matrix_reg_2__5__14_ ( .D(n3773), .CK(clk), .RN(rst_n), .QN(n435)
         );
  DFFRX1 x_matrix_reg_6__1__14_ ( .D(n4221), .CK(clk), .RN(rst_n), .QN(n579)
         );
  DFFRX1 x_matrix_reg_2__5__13_ ( .D(n3774), .CK(clk), .RN(rst_n), .QN(n436)
         );
  DFFRX1 x_matrix_reg_6__1__13_ ( .D(n4222), .CK(clk), .RN(rst_n), .QN(n580)
         );
  DFFRX1 x_matrix_reg_2__5__12_ ( .D(n3775), .CK(clk), .RN(rst_n), .QN(n437)
         );
  DFFRX1 x_matrix_reg_6__1__12_ ( .D(n4223), .CK(clk), .RN(rst_n), .QN(n581)
         );
  DFFRX1 x_matrix_reg_2__5__11_ ( .D(n3776), .CK(clk), .RN(rst_n), .QN(n438)
         );
  DFFRX1 x_matrix_reg_6__1__11_ ( .D(n4224), .CK(clk), .RN(rst_n), .QN(n582)
         );
  DFFRX1 x_matrix_reg_2__5__10_ ( .D(n3777), .CK(clk), .RN(rst_n), .QN(n439)
         );
  DFFRX1 x_matrix_reg_6__1__10_ ( .D(n4225), .CK(clk), .RN(rst_n), .QN(n583)
         );
  DFFRX1 x_matrix_reg_2__5__9_ ( .D(n3778), .CK(clk), .RN(rst_n), .QN(n440) );
  DFFRX1 x_matrix_reg_6__1__9_ ( .D(n4226), .CK(clk), .RN(rst_n), .QN(n584) );
  DFFRX1 x_matrix_reg_2__5__8_ ( .D(n3779), .CK(clk), .RN(rst_n), .QN(n441) );
  DFFRX1 x_matrix_reg_6__1__8_ ( .D(n4227), .CK(clk), .RN(rst_n), .QN(n585) );
  DFFRX1 x_matrix_reg_0__7__3_ ( .D(n3560), .CK(clk), .RN(rst_n), .QN(n382) );
  DFFRX1 x_matrix_reg_4__3__3_ ( .D(n4008), .CK(clk), .RN(rst_n), .QN(n510) );
  DFFRX1 x_matrix_reg_2__5__7_ ( .D(n3780), .CK(clk), .RN(rst_n), .QN(n442) );
  DFFRX1 x_matrix_reg_6__1__7_ ( .D(n4228), .CK(clk), .RN(rst_n), .QN(n586) );
  DFFRX1 x_matrix_reg_2__5__6_ ( .D(n3781), .CK(clk), .RN(rst_n), .QN(n443) );
  DFFRX1 x_matrix_reg_6__1__6_ ( .D(n4229), .CK(clk), .RN(rst_n), .QN(n587) );
  DFFRX1 x_matrix_reg_2__5__5_ ( .D(n3782), .CK(clk), .RN(rst_n), .QN(n444) );
  DFFRX1 x_matrix_reg_6__1__5_ ( .D(n4230), .CK(clk), .RN(rst_n), .QN(n588) );
  DFFRX1 x_matrix_reg_2__5__4_ ( .D(n3783), .CK(clk), .RN(rst_n), .QN(n445) );
  DFFRX1 x_matrix_reg_6__1__4_ ( .D(n4231), .CK(clk), .RN(rst_n), .QN(n589) );
  DFFRX1 x_matrix_reg_2__5__3_ ( .D(n3784), .CK(clk), .RN(rst_n), .QN(n446) );
  DFFRX1 x_matrix_reg_6__1__3_ ( .D(n4232), .CK(clk), .RN(rst_n), .QN(n590) );
  DFFRX1 x_matrix_reg_2__5__2_ ( .D(n3785), .CK(clk), .RN(rst_n), .QN(n447) );
  DFFRX1 x_matrix_reg_6__1__2_ ( .D(n4233), .CK(clk), .RN(rst_n), .QN(n591) );
  DFFRX1 x_matrix_reg_2__5__1_ ( .D(n3786), .CK(clk), .RN(rst_n), .QN(n448) );
  DFFRX1 x_matrix_reg_6__1__1_ ( .D(n4234), .CK(clk), .RN(rst_n), .QN(n592) );
  DFFRX1 x_matrix_reg_2__5__0_ ( .D(n3787), .CK(clk), .RN(rst_n), .QN(n449) );
  DFFRX1 x_matrix_reg_6__1__0_ ( .D(n4235), .CK(clk), .RN(rst_n), .QN(n593) );
  DFFRX1 x_matrix_reg_2__6__15_ ( .D(n3788), .CK(clk), .RN(rst_n), .QN(n450)
         );
  DFFRX1 x_matrix_reg_6__2__15_ ( .D(n4236), .CK(clk), .RN(rst_n), .QN(n594)
         );
  DFFRX1 x_matrix_reg_2__6__14_ ( .D(n3789), .CK(clk), .RN(rst_n), .QN(n451)
         );
  DFFRX1 x_matrix_reg_6__2__14_ ( .D(n4237), .CK(clk), .RN(rst_n), .QN(n595)
         );
  DFFRX1 x_matrix_reg_0__7__2_ ( .D(n3561), .CK(clk), .RN(rst_n), .QN(n383) );
  DFFRX1 x_matrix_reg_4__3__2_ ( .D(n4009), .CK(clk), .RN(rst_n), .QN(n511) );
  DFFRX1 x_matrix_reg_2__6__13_ ( .D(n3790), .CK(clk), .RN(rst_n), .QN(n452)
         );
  DFFRX1 x_matrix_reg_6__2__13_ ( .D(n4238), .CK(clk), .RN(rst_n), .QN(n596)
         );
  DFFRX1 x_matrix_reg_2__6__12_ ( .D(n3791), .CK(clk), .RN(rst_n), .QN(n453)
         );
  DFFRX1 x_matrix_reg_6__2__12_ ( .D(n4239), .CK(clk), .RN(rst_n), .QN(n597)
         );
  DFFRX1 x_matrix_reg_2__6__11_ ( .D(n3792), .CK(clk), .RN(rst_n), .QN(n454)
         );
  DFFRX1 x_matrix_reg_6__2__11_ ( .D(n4240), .CK(clk), .RN(rst_n), .QN(n598)
         );
  DFFRX1 x_matrix_reg_2__6__10_ ( .D(n3793), .CK(clk), .RN(rst_n), .QN(n455)
         );
  DFFRX1 x_matrix_reg_6__2__10_ ( .D(n4241), .CK(clk), .RN(rst_n), .QN(n599)
         );
  DFFRX1 x_matrix_reg_2__6__9_ ( .D(n3794), .CK(clk), .RN(rst_n), .QN(n456) );
  DFFRX1 x_matrix_reg_6__2__9_ ( .D(n4242), .CK(clk), .RN(rst_n), .QN(n600) );
  DFFRX1 x_matrix_reg_2__6__8_ ( .D(n3795), .CK(clk), .RN(rst_n), .QN(n457) );
  DFFRX1 x_matrix_reg_6__2__8_ ( .D(n4243), .CK(clk), .RN(rst_n), .QN(n601) );
  DFFRX1 x_matrix_reg_2__6__7_ ( .D(n3796), .CK(clk), .RN(rst_n), .QN(n458) );
  DFFRX1 x_matrix_reg_6__2__7_ ( .D(n4244), .CK(clk), .RN(rst_n), .QN(n602) );
  DFFRX1 x_matrix_reg_2__6__6_ ( .D(n3797), .CK(clk), .RN(rst_n), .QN(n459) );
  DFFRX1 x_matrix_reg_6__2__6_ ( .D(n4245), .CK(clk), .RN(rst_n), .QN(n603) );
  DFFRX1 x_matrix_reg_2__6__5_ ( .D(n3798), .CK(clk), .RN(rst_n), .QN(n460) );
  DFFRX1 x_matrix_reg_6__2__5_ ( .D(n4246), .CK(clk), .RN(rst_n), .QN(n604) );
  DFFRX1 x_matrix_reg_2__6__4_ ( .D(n3799), .CK(clk), .RN(rst_n), .QN(n461) );
  DFFRX1 x_matrix_reg_6__2__4_ ( .D(n4247), .CK(clk), .RN(rst_n), .QN(n605) );
  DFFRX1 x_matrix_reg_0__7__1_ ( .D(n3562), .CK(clk), .RN(rst_n), .QN(n384) );
  DFFRX1 x_matrix_reg_4__3__1_ ( .D(n4010), .CK(clk), .RN(rst_n), .QN(n512) );
  DFFRX1 x_matrix_reg_2__6__3_ ( .D(n3800), .CK(clk), .RN(rst_n), .QN(n462) );
  DFFRX1 x_matrix_reg_6__2__3_ ( .D(n4248), .CK(clk), .RN(rst_n), .QN(n606) );
  DFFRX1 x_matrix_reg_2__6__2_ ( .D(n3801), .CK(clk), .RN(rst_n), .QN(n463) );
  DFFRX1 x_matrix_reg_6__2__2_ ( .D(n4249), .CK(clk), .RN(rst_n), .QN(n607) );
  DFFRX1 x_matrix_reg_2__6__1_ ( .D(n3802), .CK(clk), .RN(rst_n), .QN(n464) );
  DFFRX1 x_matrix_reg_6__2__1_ ( .D(n4250), .CK(clk), .RN(rst_n), .QN(n608) );
  DFFRX1 x_matrix_reg_2__6__0_ ( .D(n3803), .CK(clk), .RN(rst_n), .QN(n465) );
  DFFRX1 x_matrix_reg_6__2__0_ ( .D(n4251), .CK(clk), .RN(rst_n), .QN(n609) );
  DFFRX1 x_matrix_reg_0__7__15_ ( .D(n3548), .CK(clk), .RN(rst_n), .QN(n370)
         );
  DFFRX1 x_matrix_reg_4__3__15_ ( .D(n3996), .CK(clk), .RN(rst_n), .QN(n498)
         );
  DFFRX1 x_matrix_reg_0__7__14_ ( .D(n3549), .CK(clk), .RN(rst_n), .QN(n371)
         );
  DFFRX1 x_matrix_reg_4__3__14_ ( .D(n3997), .CK(clk), .RN(rst_n), .QN(n499)
         );
  DFFRX1 x_matrix_reg_0__7__13_ ( .D(n3550), .CK(clk), .RN(rst_n), .QN(n372)
         );
  DFFRX1 x_matrix_reg_4__3__13_ ( .D(n3998), .CK(clk), .RN(rst_n), .QN(n500)
         );
  DFFRX1 x_matrix_reg_0__7__12_ ( .D(n3551), .CK(clk), .RN(rst_n), .QN(n373)
         );
  DFFRX1 x_matrix_reg_4__3__12_ ( .D(n3999), .CK(clk), .RN(rst_n), .QN(n501)
         );
  DFFRX1 x_matrix_reg_0__7__11_ ( .D(n3552), .CK(clk), .RN(rst_n), .QN(n374)
         );
  DFFRX1 x_matrix_reg_4__3__11_ ( .D(n4000), .CK(clk), .RN(rst_n), .QN(n502)
         );
  DFFRX1 x_matrix_reg_0__7__10_ ( .D(n3553), .CK(clk), .RN(rst_n), .QN(n375)
         );
  DFFRX1 x_matrix_reg_4__3__10_ ( .D(n4001), .CK(clk), .RN(rst_n), .QN(n503)
         );
  DFFRX1 x_matrix_reg_0__7__0_ ( .D(n3563), .CK(clk), .RN(rst_n), .QN(n385) );
  DFFRX1 x_matrix_reg_4__3__0_ ( .D(n4011), .CK(clk), .RN(rst_n), .QN(n513) );
  DFFSX1 in_addr_cnt_reg_9_ ( .D(n4460), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[9]), .QN(n4496) );
  DFFRHQX1 x_matrix_reg_0__3__9_ ( .D(n3490), .CK(clk), .RN(rst_n), .Q(
        x_matrix[713]) );
  DFFRHQX1 x_matrix_reg_2__3__9_ ( .D(n3746), .CK(clk), .RN(rst_n), .Q(
        x_matrix[489]) );
  DFFRHQX1 x_matrix_reg_4__7__9_ ( .D(n4066), .CK(clk), .RN(rst_n), .Q(
        x_matrix[265]) );
  DFFRHQX1 x_matrix_reg_6__7__9_ ( .D(n4322), .CK(clk), .RN(rst_n), .Q(
        x_matrix[89]) );
  DFFRHQX1 x_matrix_reg_0__3__8_ ( .D(n3491), .CK(clk), .RN(rst_n), .Q(
        x_matrix[712]) );
  DFFRHQX1 x_matrix_reg_2__3__8_ ( .D(n3747), .CK(clk), .RN(rst_n), .Q(
        x_matrix[488]) );
  DFFRHQX1 x_matrix_reg_4__7__8_ ( .D(n4067), .CK(clk), .RN(rst_n), .Q(
        x_matrix[264]) );
  DFFRHQX1 x_matrix_reg_6__7__8_ ( .D(n4323), .CK(clk), .RN(rst_n), .Q(
        x_matrix[88]) );
  DFFRHQX1 x_matrix_reg_0__3__7_ ( .D(n3492), .CK(clk), .RN(rst_n), .Q(
        x_matrix[711]) );
  DFFRHQX1 x_matrix_reg_2__3__7_ ( .D(n3748), .CK(clk), .RN(rst_n), .Q(
        x_matrix[487]) );
  DFFRHQX1 x_matrix_reg_4__7__7_ ( .D(n4068), .CK(clk), .RN(rst_n), .Q(
        x_matrix[263]) );
  DFFRHQX1 x_matrix_reg_6__7__7_ ( .D(n4324), .CK(clk), .RN(rst_n), .Q(
        x_matrix[87]) );
  DFFRHQX1 x_matrix_reg_0__3__6_ ( .D(n3493), .CK(clk), .RN(rst_n), .Q(
        x_matrix[710]) );
  DFFRHQX1 x_matrix_reg_2__3__6_ ( .D(n3749), .CK(clk), .RN(rst_n), .Q(
        x_matrix[486]) );
  DFFRHQX1 x_matrix_reg_4__7__6_ ( .D(n4069), .CK(clk), .RN(rst_n), .Q(
        x_matrix[262]) );
  DFFRHQX1 x_matrix_reg_6__7__6_ ( .D(n4325), .CK(clk), .RN(rst_n), .Q(
        x_matrix[86]) );
  DFFRHQX1 x_matrix_reg_0__0__15_ ( .D(n3436), .CK(clk), .RN(rst_n), .Q(
        x_matrix[767]) );
  DFFRHQX1 x_matrix_reg_0__4__15_ ( .D(n3500), .CK(clk), .RN(rst_n), .Q(
        x_matrix[703]) );
  DFFRHQX1 x_matrix_reg_2__0__15_ ( .D(n3692), .CK(clk), .RN(rst_n), .Q(
        x_matrix[543]) );
  DFFRHQX1 x_matrix_reg_2__4__15_ ( .D(n3756), .CK(clk), .RN(rst_n), .Q(
        x_matrix[479]) );
  DFFRHQX1 x_matrix_reg_0__0__14_ ( .D(n3437), .CK(clk), .RN(rst_n), .Q(
        x_matrix[766]) );
  DFFRHQX1 x_matrix_reg_0__4__14_ ( .D(n3501), .CK(clk), .RN(rst_n), .Q(
        x_matrix[702]) );
  DFFRHQX1 x_matrix_reg_2__0__14_ ( .D(n3693), .CK(clk), .RN(rst_n), .Q(
        x_matrix[542]) );
  DFFRHQX1 x_matrix_reg_2__4__14_ ( .D(n3757), .CK(clk), .RN(rst_n), .Q(
        x_matrix[478]) );
  DFFRHQX1 x_matrix_reg_0__0__13_ ( .D(n3438), .CK(clk), .RN(rst_n), .Q(
        x_matrix[765]) );
  DFFRHQX1 x_matrix_reg_0__4__13_ ( .D(n3502), .CK(clk), .RN(rst_n), .Q(
        x_matrix[701]) );
  DFFRHQX1 x_matrix_reg_2__0__13_ ( .D(n3694), .CK(clk), .RN(rst_n), .Q(
        x_matrix[541]) );
  DFFRHQX1 x_matrix_reg_2__4__13_ ( .D(n3758), .CK(clk), .RN(rst_n), .Q(
        x_matrix[477]) );
  DFFRHQX1 x_matrix_reg_0__0__12_ ( .D(n3439), .CK(clk), .RN(rst_n), .Q(
        x_matrix[764]) );
  DFFRHQX1 x_matrix_reg_0__4__12_ ( .D(n3503), .CK(clk), .RN(rst_n), .Q(
        x_matrix[700]) );
  DFFRHQX1 x_matrix_reg_2__0__12_ ( .D(n3695), .CK(clk), .RN(rst_n), .Q(
        x_matrix[540]) );
  DFFRHQX1 x_matrix_reg_2__4__12_ ( .D(n3759), .CK(clk), .RN(rst_n), .Q(
        x_matrix[476]) );
  DFFRHQX1 x_matrix_reg_0__3__5_ ( .D(n3494), .CK(clk), .RN(rst_n), .Q(
        x_matrix[709]) );
  DFFRHQX1 x_matrix_reg_2__3__5_ ( .D(n3750), .CK(clk), .RN(rst_n), .Q(
        x_matrix[485]) );
  DFFRHQX1 x_matrix_reg_4__7__5_ ( .D(n4070), .CK(clk), .RN(rst_n), .Q(
        x_matrix[261]) );
  DFFRHQX1 x_matrix_reg_6__7__5_ ( .D(n4326), .CK(clk), .RN(rst_n), .Q(
        x_matrix[85]) );
  DFFRHQX1 x_matrix_reg_0__0__11_ ( .D(n3440), .CK(clk), .RN(rst_n), .Q(
        x_matrix[763]) );
  DFFRHQX1 x_matrix_reg_0__4__11_ ( .D(n3504), .CK(clk), .RN(rst_n), .Q(
        x_matrix[699]) );
  DFFRHQX1 x_matrix_reg_2__0__11_ ( .D(n3696), .CK(clk), .RN(rst_n), .Q(
        x_matrix[539]) );
  DFFRHQX1 x_matrix_reg_2__4__11_ ( .D(n3760), .CK(clk), .RN(rst_n), .Q(
        x_matrix[475]) );
  DFFRHQX1 x_matrix_reg_0__0__10_ ( .D(n3441), .CK(clk), .RN(rst_n), .Q(
        x_matrix[762]) );
  DFFRHQX1 x_matrix_reg_0__4__10_ ( .D(n3505), .CK(clk), .RN(rst_n), .Q(
        x_matrix[698]) );
  DFFRHQX1 x_matrix_reg_2__0__10_ ( .D(n3697), .CK(clk), .RN(rst_n), .Q(
        x_matrix[538]) );
  DFFRHQX1 x_matrix_reg_2__4__10_ ( .D(n3761), .CK(clk), .RN(rst_n), .Q(
        x_matrix[474]) );
  DFFRHQX1 x_matrix_reg_0__0__9_ ( .D(n3442), .CK(clk), .RN(rst_n), .Q(
        x_matrix[761]) );
  DFFRHQX1 x_matrix_reg_0__4__9_ ( .D(n3506), .CK(clk), .RN(rst_n), .Q(
        x_matrix[697]) );
  DFFRHQX1 x_matrix_reg_2__0__9_ ( .D(n3698), .CK(clk), .RN(rst_n), .Q(
        x_matrix[537]) );
  DFFRHQX1 x_matrix_reg_2__4__9_ ( .D(n3762), .CK(clk), .RN(rst_n), .Q(
        x_matrix[473]) );
  DFFRHQX1 x_matrix_reg_0__0__8_ ( .D(n3443), .CK(clk), .RN(rst_n), .Q(
        x_matrix[760]) );
  DFFRHQX1 x_matrix_reg_0__4__8_ ( .D(n3507), .CK(clk), .RN(rst_n), .Q(
        x_matrix[696]) );
  DFFRHQX1 x_matrix_reg_2__0__8_ ( .D(n3699), .CK(clk), .RN(rst_n), .Q(
        x_matrix[536]) );
  DFFRHQX1 x_matrix_reg_2__4__8_ ( .D(n3763), .CK(clk), .RN(rst_n), .Q(
        x_matrix[472]) );
  DFFRHQX1 x_matrix_reg_0__0__7_ ( .D(n3444), .CK(clk), .RN(rst_n), .Q(
        x_matrix[759]) );
  DFFRHQX1 x_matrix_reg_0__4__7_ ( .D(n3508), .CK(clk), .RN(rst_n), .Q(
        x_matrix[695]) );
  DFFRHQX1 x_matrix_reg_2__0__7_ ( .D(n3700), .CK(clk), .RN(rst_n), .Q(
        x_matrix[535]) );
  DFFRHQX1 x_matrix_reg_2__4__7_ ( .D(n3764), .CK(clk), .RN(rst_n), .Q(
        x_matrix[471]) );
  DFFRHQX1 x_matrix_reg_0__0__6_ ( .D(n3445), .CK(clk), .RN(rst_n), .Q(
        x_matrix[758]) );
  DFFRHQX1 x_matrix_reg_0__4__6_ ( .D(n3509), .CK(clk), .RN(rst_n), .Q(
        x_matrix[694]) );
  DFFRHQX1 x_matrix_reg_2__0__6_ ( .D(n3701), .CK(clk), .RN(rst_n), .Q(
        x_matrix[534]) );
  DFFRHQX1 x_matrix_reg_2__4__6_ ( .D(n3765), .CK(clk), .RN(rst_n), .Q(
        x_matrix[470]) );
  DFFRHQX1 x_matrix_reg_0__0__5_ ( .D(n3446), .CK(clk), .RN(rst_n), .Q(
        x_matrix[757]) );
  DFFRHQX1 x_matrix_reg_0__4__5_ ( .D(n3510), .CK(clk), .RN(rst_n), .Q(
        x_matrix[693]) );
  DFFRHQX1 x_matrix_reg_2__0__5_ ( .D(n3702), .CK(clk), .RN(rst_n), .Q(
        x_matrix[533]) );
  DFFRHQX1 x_matrix_reg_2__4__5_ ( .D(n3766), .CK(clk), .RN(rst_n), .Q(
        x_matrix[469]) );
  DFFRHQX1 x_matrix_reg_0__0__4_ ( .D(n3447), .CK(clk), .RN(rst_n), .Q(
        x_matrix[756]) );
  DFFRHQX1 x_matrix_reg_0__4__4_ ( .D(n3511), .CK(clk), .RN(rst_n), .Q(
        x_matrix[692]) );
  DFFRHQX1 x_matrix_reg_2__0__4_ ( .D(n3703), .CK(clk), .RN(rst_n), .Q(
        x_matrix[532]) );
  DFFRHQX1 x_matrix_reg_2__4__4_ ( .D(n3767), .CK(clk), .RN(rst_n), .Q(
        x_matrix[468]) );
  DFFRHQX1 x_matrix_reg_0__0__3_ ( .D(n3448), .CK(clk), .RN(rst_n), .Q(
        x_matrix[755]) );
  DFFRHQX1 x_matrix_reg_0__4__3_ ( .D(n3512), .CK(clk), .RN(rst_n), .Q(
        x_matrix[691]) );
  DFFRHQX1 x_matrix_reg_2__0__3_ ( .D(n3704), .CK(clk), .RN(rst_n), .Q(
        x_matrix[531]) );
  DFFRHQX1 x_matrix_reg_2__4__3_ ( .D(n3768), .CK(clk), .RN(rst_n), .Q(
        x_matrix[467]) );
  DFFRHQX1 x_matrix_reg_0__0__2_ ( .D(n3449), .CK(clk), .RN(rst_n), .Q(
        x_matrix[754]) );
  DFFRHQX1 x_matrix_reg_0__4__2_ ( .D(n3513), .CK(clk), .RN(rst_n), .Q(
        x_matrix[690]) );
  DFFRHQX1 x_matrix_reg_2__0__2_ ( .D(n3705), .CK(clk), .RN(rst_n), .Q(
        x_matrix[530]) );
  DFFRHQX1 x_matrix_reg_2__4__2_ ( .D(n3769), .CK(clk), .RN(rst_n), .Q(
        x_matrix[466]) );
  DFFRHQX1 x_matrix_reg_0__3__4_ ( .D(n3495), .CK(clk), .RN(rst_n), .Q(
        x_matrix[708]) );
  DFFRHQX1 x_matrix_reg_2__3__4_ ( .D(n3751), .CK(clk), .RN(rst_n), .Q(
        x_matrix[484]) );
  DFFRHQX1 x_matrix_reg_4__7__4_ ( .D(n4071), .CK(clk), .RN(rst_n), .Q(
        x_matrix[260]) );
  DFFRHQX1 x_matrix_reg_6__7__4_ ( .D(n4327), .CK(clk), .RN(rst_n), .Q(
        x_matrix[84]) );
  DFFRHQX1 x_matrix_reg_0__0__1_ ( .D(n3450), .CK(clk), .RN(rst_n), .Q(
        x_matrix[753]) );
  DFFRHQX1 x_matrix_reg_0__4__1_ ( .D(n3514), .CK(clk), .RN(rst_n), .Q(
        x_matrix[689]) );
  DFFRHQX1 x_matrix_reg_2__0__1_ ( .D(n3706), .CK(clk), .RN(rst_n), .Q(
        x_matrix[529]) );
  DFFRHQX1 x_matrix_reg_2__4__1_ ( .D(n3770), .CK(clk), .RN(rst_n), .Q(
        x_matrix[465]) );
  DFFRHQX1 x_matrix_reg_0__0__0_ ( .D(n3451), .CK(clk), .RN(rst_n), .Q(
        x_matrix[752]) );
  DFFRHQX1 x_matrix_reg_0__4__0_ ( .D(n3515), .CK(clk), .RN(rst_n), .Q(
        x_matrix[688]) );
  DFFRHQX1 x_matrix_reg_2__0__0_ ( .D(n3707), .CK(clk), .RN(rst_n), .Q(
        x_matrix[528]) );
  DFFRHQX1 x_matrix_reg_2__4__0_ ( .D(n3771), .CK(clk), .RN(rst_n), .Q(
        x_matrix[464]) );
  DFFRHQX1 x_matrix_reg_0__1__15_ ( .D(n3452), .CK(clk), .RN(rst_n), .Q(
        x_matrix[751]) );
  DFFRHQX1 x_matrix_reg_2__1__15_ ( .D(n3708), .CK(clk), .RN(rst_n), .Q(
        x_matrix[527]) );
  DFFRHQX1 x_matrix_reg_4__5__15_ ( .D(n4028), .CK(clk), .RN(rst_n), .Q(
        x_matrix[303]) );
  DFFRHQX1 x_matrix_reg_6__5__15_ ( .D(n4284), .CK(clk), .RN(rst_n), .Q(
        x_matrix[127]) );
  DFFRHQX1 x_matrix_reg_0__1__14_ ( .D(n3453), .CK(clk), .RN(rst_n), .Q(
        x_matrix[750]) );
  DFFRHQX1 x_matrix_reg_2__1__14_ ( .D(n3709), .CK(clk), .RN(rst_n), .Q(
        x_matrix[526]) );
  DFFRHQX1 x_matrix_reg_4__5__14_ ( .D(n4029), .CK(clk), .RN(rst_n), .Q(
        x_matrix[302]) );
  DFFRHQX1 x_matrix_reg_6__5__14_ ( .D(n4285), .CK(clk), .RN(rst_n), .Q(
        x_matrix[126]) );
  DFFRHQX1 x_matrix_reg_0__1__13_ ( .D(n3454), .CK(clk), .RN(rst_n), .Q(
        x_matrix[749]) );
  DFFRHQX1 x_matrix_reg_2__1__13_ ( .D(n3710), .CK(clk), .RN(rst_n), .Q(
        x_matrix[525]) );
  DFFRHQX1 x_matrix_reg_4__5__13_ ( .D(n4030), .CK(clk), .RN(rst_n), .Q(
        x_matrix[301]) );
  DFFRHQX1 x_matrix_reg_6__5__13_ ( .D(n4286), .CK(clk), .RN(rst_n), .Q(
        x_matrix[125]) );
  DFFRHQX1 x_matrix_reg_0__1__12_ ( .D(n3455), .CK(clk), .RN(rst_n), .Q(
        x_matrix[748]) );
  DFFRHQX1 x_matrix_reg_2__1__12_ ( .D(n3711), .CK(clk), .RN(rst_n), .Q(
        x_matrix[524]) );
  DFFRHQX1 x_matrix_reg_4__5__12_ ( .D(n4031), .CK(clk), .RN(rst_n), .Q(
        x_matrix[300]) );
  DFFRHQX1 x_matrix_reg_6__5__12_ ( .D(n4287), .CK(clk), .RN(rst_n), .Q(
        x_matrix[124]) );
  DFFRHQX1 x_matrix_reg_0__1__11_ ( .D(n3456), .CK(clk), .RN(rst_n), .Q(
        x_matrix[747]) );
  DFFRHQX1 x_matrix_reg_2__1__11_ ( .D(n3712), .CK(clk), .RN(rst_n), .Q(
        x_matrix[523]) );
  DFFRHQX1 x_matrix_reg_4__5__11_ ( .D(n4032), .CK(clk), .RN(rst_n), .Q(
        x_matrix[299]) );
  DFFRHQX1 x_matrix_reg_6__5__11_ ( .D(n4288), .CK(clk), .RN(rst_n), .Q(
        x_matrix[123]) );
  DFFRHQX1 x_matrix_reg_0__1__10_ ( .D(n3457), .CK(clk), .RN(rst_n), .Q(
        x_matrix[746]) );
  DFFRHQX1 x_matrix_reg_2__1__10_ ( .D(n3713), .CK(clk), .RN(rst_n), .Q(
        x_matrix[522]) );
  DFFRHQX1 x_matrix_reg_4__5__10_ ( .D(n4033), .CK(clk), .RN(rst_n), .Q(
        x_matrix[298]) );
  DFFRHQX1 x_matrix_reg_6__5__10_ ( .D(n4289), .CK(clk), .RN(rst_n), .Q(
        x_matrix[122]) );
  DFFRHQX1 x_matrix_reg_0__1__9_ ( .D(n3458), .CK(clk), .RN(rst_n), .Q(
        x_matrix[745]) );
  DFFRHQX1 x_matrix_reg_2__1__9_ ( .D(n3714), .CK(clk), .RN(rst_n), .Q(
        x_matrix[521]) );
  DFFRHQX1 x_matrix_reg_4__5__9_ ( .D(n4034), .CK(clk), .RN(rst_n), .Q(
        x_matrix[297]) );
  DFFRHQX1 x_matrix_reg_6__5__9_ ( .D(n4290), .CK(clk), .RN(rst_n), .Q(
        x_matrix[121]) );
  DFFRHQX1 x_matrix_reg_0__1__8_ ( .D(n3459), .CK(clk), .RN(rst_n), .Q(
        x_matrix[744]) );
  DFFRHQX1 x_matrix_reg_2__1__8_ ( .D(n3715), .CK(clk), .RN(rst_n), .Q(
        x_matrix[520]) );
  DFFRHQX1 x_matrix_reg_4__5__8_ ( .D(n4035), .CK(clk), .RN(rst_n), .Q(
        x_matrix[296]) );
  DFFRHQX1 x_matrix_reg_6__5__8_ ( .D(n4291), .CK(clk), .RN(rst_n), .Q(
        x_matrix[120]) );
  DFFRHQX1 x_matrix_reg_0__3__3_ ( .D(n3496), .CK(clk), .RN(rst_n), .Q(
        x_matrix[707]) );
  DFFRHQX1 x_matrix_reg_2__3__3_ ( .D(n3752), .CK(clk), .RN(rst_n), .Q(
        x_matrix[483]) );
  DFFRHQX1 x_matrix_reg_4__7__3_ ( .D(n4072), .CK(clk), .RN(rst_n), .Q(
        x_matrix[259]) );
  DFFRHQX1 x_matrix_reg_6__7__3_ ( .D(n4328), .CK(clk), .RN(rst_n), .Q(
        x_matrix[83]) );
  DFFRHQX1 x_matrix_reg_0__1__7_ ( .D(n3460), .CK(clk), .RN(rst_n), .Q(
        x_matrix[743]) );
  DFFRHQX1 x_matrix_reg_2__1__7_ ( .D(n3716), .CK(clk), .RN(rst_n), .Q(
        x_matrix[519]) );
  DFFRHQX1 x_matrix_reg_4__5__7_ ( .D(n4036), .CK(clk), .RN(rst_n), .Q(
        x_matrix[295]) );
  DFFRHQX1 x_matrix_reg_6__5__7_ ( .D(n4292), .CK(clk), .RN(rst_n), .Q(
        x_matrix[119]) );
  DFFRHQX1 x_matrix_reg_0__1__6_ ( .D(n3461), .CK(clk), .RN(rst_n), .Q(
        x_matrix[742]) );
  DFFRHQX1 x_matrix_reg_2__1__6_ ( .D(n3717), .CK(clk), .RN(rst_n), .Q(
        x_matrix[518]) );
  DFFRHQX1 x_matrix_reg_4__5__6_ ( .D(n4037), .CK(clk), .RN(rst_n), .Q(
        x_matrix[294]) );
  DFFRHQX1 x_matrix_reg_6__5__6_ ( .D(n4293), .CK(clk), .RN(rst_n), .Q(
        x_matrix[118]) );
  DFFRHQX1 x_matrix_reg_0__1__5_ ( .D(n3462), .CK(clk), .RN(rst_n), .Q(
        x_matrix[741]) );
  DFFRHQX1 x_matrix_reg_2__1__5_ ( .D(n3718), .CK(clk), .RN(rst_n), .Q(
        x_matrix[517]) );
  DFFRHQX1 x_matrix_reg_4__5__5_ ( .D(n4038), .CK(clk), .RN(rst_n), .Q(
        x_matrix[293]) );
  DFFRHQX1 x_matrix_reg_6__5__5_ ( .D(n4294), .CK(clk), .RN(rst_n), .Q(
        x_matrix[117]) );
  DFFRHQX1 x_matrix_reg_0__1__4_ ( .D(n3463), .CK(clk), .RN(rst_n), .Q(
        x_matrix[740]) );
  DFFRHQX1 x_matrix_reg_2__1__4_ ( .D(n3719), .CK(clk), .RN(rst_n), .Q(
        x_matrix[516]) );
  DFFRHQX1 x_matrix_reg_4__5__4_ ( .D(n4039), .CK(clk), .RN(rst_n), .Q(
        x_matrix[292]) );
  DFFRHQX1 x_matrix_reg_6__5__4_ ( .D(n4295), .CK(clk), .RN(rst_n), .Q(
        x_matrix[116]) );
  DFFRHQX1 x_matrix_reg_0__1__3_ ( .D(n3464), .CK(clk), .RN(rst_n), .Q(
        x_matrix[739]) );
  DFFRHQX1 x_matrix_reg_2__1__3_ ( .D(n3720), .CK(clk), .RN(rst_n), .Q(
        x_matrix[515]) );
  DFFRHQX1 x_matrix_reg_4__5__3_ ( .D(n4040), .CK(clk), .RN(rst_n), .Q(
        x_matrix[291]) );
  DFFRHQX1 x_matrix_reg_6__5__3_ ( .D(n4296), .CK(clk), .RN(rst_n), .Q(
        x_matrix[115]) );
  DFFRHQX1 x_matrix_reg_0__1__2_ ( .D(n3465), .CK(clk), .RN(rst_n), .Q(
        x_matrix[738]) );
  DFFRHQX1 x_matrix_reg_2__1__2_ ( .D(n3721), .CK(clk), .RN(rst_n), .Q(
        x_matrix[514]) );
  DFFRHQX1 x_matrix_reg_4__5__2_ ( .D(n4041), .CK(clk), .RN(rst_n), .Q(
        x_matrix[290]) );
  DFFRHQX1 x_matrix_reg_6__5__2_ ( .D(n4297), .CK(clk), .RN(rst_n), .Q(
        x_matrix[114]) );
  DFFRHQX1 x_matrix_reg_0__1__1_ ( .D(n3466), .CK(clk), .RN(rst_n), .Q(
        x_matrix[737]) );
  DFFRHQX1 x_matrix_reg_2__1__1_ ( .D(n3722), .CK(clk), .RN(rst_n), .Q(
        x_matrix[513]) );
  DFFRHQX1 x_matrix_reg_4__5__1_ ( .D(n4042), .CK(clk), .RN(rst_n), .Q(
        x_matrix[289]) );
  DFFRHQX1 x_matrix_reg_6__5__1_ ( .D(n4298), .CK(clk), .RN(rst_n), .Q(
        x_matrix[113]) );
  DFFRHQX1 x_matrix_reg_0__1__0_ ( .D(n3467), .CK(clk), .RN(rst_n), .Q(
        x_matrix[736]) );
  DFFRHQX1 x_matrix_reg_2__1__0_ ( .D(n3723), .CK(clk), .RN(rst_n), .Q(
        x_matrix[512]) );
  DFFRHQX1 x_matrix_reg_4__5__0_ ( .D(n4043), .CK(clk), .RN(rst_n), .Q(
        x_matrix[288]) );
  DFFRHQX1 x_matrix_reg_6__5__0_ ( .D(n4299), .CK(clk), .RN(rst_n), .Q(
        x_matrix[112]) );
  DFFRHQX1 x_matrix_reg_0__2__15_ ( .D(n3468), .CK(clk), .RN(rst_n), .Q(
        x_matrix[735]) );
  DFFRHQX1 x_matrix_reg_2__2__15_ ( .D(n3724), .CK(clk), .RN(rst_n), .Q(
        x_matrix[511]) );
  DFFRHQX1 x_matrix_reg_4__6__15_ ( .D(n4044), .CK(clk), .RN(rst_n), .Q(
        x_matrix[287]) );
  DFFRHQX1 x_matrix_reg_6__6__15_ ( .D(n4300), .CK(clk), .RN(rst_n), .Q(
        x_matrix[111]) );
  DFFRHQX1 x_matrix_reg_0__2__14_ ( .D(n3469), .CK(clk), .RN(rst_n), .Q(
        x_matrix[734]) );
  DFFRHQX1 x_matrix_reg_2__2__14_ ( .D(n3725), .CK(clk), .RN(rst_n), .Q(
        x_matrix[510]) );
  DFFRHQX1 x_matrix_reg_4__6__14_ ( .D(n4045), .CK(clk), .RN(rst_n), .Q(
        x_matrix[286]) );
  DFFRHQX1 x_matrix_reg_6__6__14_ ( .D(n4301), .CK(clk), .RN(rst_n), .Q(
        x_matrix[110]) );
  DFFRHQX1 x_matrix_reg_0__3__2_ ( .D(n3497), .CK(clk), .RN(rst_n), .Q(
        x_matrix[706]) );
  DFFRHQX1 x_matrix_reg_2__3__2_ ( .D(n3753), .CK(clk), .RN(rst_n), .Q(
        x_matrix[482]) );
  DFFRHQX1 x_matrix_reg_4__7__2_ ( .D(n4073), .CK(clk), .RN(rst_n), .Q(
        x_matrix[258]) );
  DFFRHQX1 x_matrix_reg_6__7__2_ ( .D(n4329), .CK(clk), .RN(rst_n), .Q(
        x_matrix[82]) );
  DFFRHQX1 x_matrix_reg_0__2__13_ ( .D(n3470), .CK(clk), .RN(rst_n), .Q(
        x_matrix[733]) );
  DFFRHQX1 x_matrix_reg_2__2__13_ ( .D(n3726), .CK(clk), .RN(rst_n), .Q(
        x_matrix[509]) );
  DFFRHQX1 x_matrix_reg_4__6__13_ ( .D(n4046), .CK(clk), .RN(rst_n), .Q(
        x_matrix[285]) );
  DFFRHQX1 x_matrix_reg_6__6__13_ ( .D(n4302), .CK(clk), .RN(rst_n), .Q(
        x_matrix[109]) );
  DFFRHQX1 x_matrix_reg_0__2__12_ ( .D(n3471), .CK(clk), .RN(rst_n), .Q(
        x_matrix[732]) );
  DFFRHQX1 x_matrix_reg_2__2__12_ ( .D(n3727), .CK(clk), .RN(rst_n), .Q(
        x_matrix[508]) );
  DFFRHQX1 x_matrix_reg_4__6__12_ ( .D(n4047), .CK(clk), .RN(rst_n), .Q(
        x_matrix[284]) );
  DFFRHQX1 x_matrix_reg_6__6__12_ ( .D(n4303), .CK(clk), .RN(rst_n), .Q(
        x_matrix[108]) );
  DFFRHQX1 x_matrix_reg_0__2__11_ ( .D(n3472), .CK(clk), .RN(rst_n), .Q(
        x_matrix[731]) );
  DFFRHQX1 x_matrix_reg_2__2__11_ ( .D(n3728), .CK(clk), .RN(rst_n), .Q(
        x_matrix[507]) );
  DFFRHQX1 x_matrix_reg_4__6__11_ ( .D(n4048), .CK(clk), .RN(rst_n), .Q(
        x_matrix[283]) );
  DFFRHQX1 x_matrix_reg_6__6__11_ ( .D(n4304), .CK(clk), .RN(rst_n), .Q(
        x_matrix[107]) );
  DFFRHQX1 x_matrix_reg_0__2__10_ ( .D(n3473), .CK(clk), .RN(rst_n), .Q(
        x_matrix[730]) );
  DFFRHQX1 x_matrix_reg_2__2__10_ ( .D(n3729), .CK(clk), .RN(rst_n), .Q(
        x_matrix[506]) );
  DFFRHQX1 x_matrix_reg_4__6__10_ ( .D(n4049), .CK(clk), .RN(rst_n), .Q(
        x_matrix[282]) );
  DFFRHQX1 x_matrix_reg_6__6__10_ ( .D(n4305), .CK(clk), .RN(rst_n), .Q(
        x_matrix[106]) );
  DFFRHQX1 x_matrix_reg_0__2__9_ ( .D(n3474), .CK(clk), .RN(rst_n), .Q(
        x_matrix[729]) );
  DFFRHQX1 x_matrix_reg_2__2__9_ ( .D(n3730), .CK(clk), .RN(rst_n), .Q(
        x_matrix[505]) );
  DFFRHQX1 x_matrix_reg_4__6__9_ ( .D(n4050), .CK(clk), .RN(rst_n), .Q(
        x_matrix[281]) );
  DFFRHQX1 x_matrix_reg_6__6__9_ ( .D(n4306), .CK(clk), .RN(rst_n), .Q(
        x_matrix[105]) );
  DFFRHQX1 x_matrix_reg_0__2__8_ ( .D(n3475), .CK(clk), .RN(rst_n), .Q(
        x_matrix[728]) );
  DFFRHQX1 x_matrix_reg_2__2__8_ ( .D(n3731), .CK(clk), .RN(rst_n), .Q(
        x_matrix[504]) );
  DFFRHQX1 x_matrix_reg_4__6__8_ ( .D(n4051), .CK(clk), .RN(rst_n), .Q(
        x_matrix[280]) );
  DFFRHQX1 x_matrix_reg_6__6__8_ ( .D(n4307), .CK(clk), .RN(rst_n), .Q(
        x_matrix[104]) );
  DFFRHQX1 x_matrix_reg_0__2__7_ ( .D(n3476), .CK(clk), .RN(rst_n), .Q(
        x_matrix[727]) );
  DFFRHQX1 x_matrix_reg_2__2__7_ ( .D(n3732), .CK(clk), .RN(rst_n), .Q(
        x_matrix[503]) );
  DFFRHQX1 x_matrix_reg_4__6__7_ ( .D(n4052), .CK(clk), .RN(rst_n), .Q(
        x_matrix[279]) );
  DFFRHQX1 x_matrix_reg_6__6__7_ ( .D(n4308), .CK(clk), .RN(rst_n), .Q(
        x_matrix[103]) );
  DFFRHQX1 x_matrix_reg_0__2__6_ ( .D(n3477), .CK(clk), .RN(rst_n), .Q(
        x_matrix[726]) );
  DFFRHQX1 x_matrix_reg_2__2__6_ ( .D(n3733), .CK(clk), .RN(rst_n), .Q(
        x_matrix[502]) );
  DFFRHQX1 x_matrix_reg_4__6__6_ ( .D(n4053), .CK(clk), .RN(rst_n), .Q(
        x_matrix[278]) );
  DFFRHQX1 x_matrix_reg_6__6__6_ ( .D(n4309), .CK(clk), .RN(rst_n), .Q(
        x_matrix[102]) );
  DFFRHQX1 x_matrix_reg_0__2__5_ ( .D(n3478), .CK(clk), .RN(rst_n), .Q(
        x_matrix[725]) );
  DFFRHQX1 x_matrix_reg_2__2__5_ ( .D(n3734), .CK(clk), .RN(rst_n), .Q(
        x_matrix[501]) );
  DFFRHQX1 x_matrix_reg_4__6__5_ ( .D(n4054), .CK(clk), .RN(rst_n), .Q(
        x_matrix[277]) );
  DFFRHQX1 x_matrix_reg_6__6__5_ ( .D(n4310), .CK(clk), .RN(rst_n), .Q(
        x_matrix[101]) );
  DFFRHQX1 x_matrix_reg_0__2__4_ ( .D(n3479), .CK(clk), .RN(rst_n), .Q(
        x_matrix[724]) );
  DFFRHQX1 x_matrix_reg_2__2__4_ ( .D(n3735), .CK(clk), .RN(rst_n), .Q(
        x_matrix[500]) );
  DFFRHQX1 x_matrix_reg_4__6__4_ ( .D(n4055), .CK(clk), .RN(rst_n), .Q(
        x_matrix[276]) );
  DFFRHQX1 x_matrix_reg_6__6__4_ ( .D(n4311), .CK(clk), .RN(rst_n), .Q(
        x_matrix[100]) );
  DFFRHQX1 x_matrix_reg_0__3__1_ ( .D(n3498), .CK(clk), .RN(rst_n), .Q(
        x_matrix[705]) );
  DFFRHQX1 x_matrix_reg_2__3__1_ ( .D(n3754), .CK(clk), .RN(rst_n), .Q(
        x_matrix[481]) );
  DFFRHQX1 x_matrix_reg_4__7__1_ ( .D(n4074), .CK(clk), .RN(rst_n), .Q(
        x_matrix[257]) );
  DFFRHQX1 x_matrix_reg_6__7__1_ ( .D(n4330), .CK(clk), .RN(rst_n), .Q(
        x_matrix[81]) );
  DFFRHQX1 x_matrix_reg_0__2__3_ ( .D(n3480), .CK(clk), .RN(rst_n), .Q(
        x_matrix[723]) );
  DFFRHQX1 x_matrix_reg_2__2__3_ ( .D(n3736), .CK(clk), .RN(rst_n), .Q(
        x_matrix[499]) );
  DFFRHQX1 x_matrix_reg_4__6__3_ ( .D(n4056), .CK(clk), .RN(rst_n), .Q(
        x_matrix[275]) );
  DFFRHQX1 x_matrix_reg_6__6__3_ ( .D(n4312), .CK(clk), .RN(rst_n), .Q(
        x_matrix[99]) );
  DFFRHQX1 x_matrix_reg_0__2__2_ ( .D(n3481), .CK(clk), .RN(rst_n), .Q(
        x_matrix[722]) );
  DFFRHQX1 x_matrix_reg_2__2__2_ ( .D(n3737), .CK(clk), .RN(rst_n), .Q(
        x_matrix[498]) );
  DFFRHQX1 x_matrix_reg_4__6__2_ ( .D(n4057), .CK(clk), .RN(rst_n), .Q(
        x_matrix[274]) );
  DFFRHQX1 x_matrix_reg_6__6__2_ ( .D(n4313), .CK(clk), .RN(rst_n), .Q(
        x_matrix[98]) );
  DFFRHQX1 x_matrix_reg_0__2__1_ ( .D(n3482), .CK(clk), .RN(rst_n), .Q(
        x_matrix[721]) );
  DFFRHQX1 x_matrix_reg_2__2__1_ ( .D(n3738), .CK(clk), .RN(rst_n), .Q(
        x_matrix[497]) );
  DFFRHQX1 x_matrix_reg_4__6__1_ ( .D(n4058), .CK(clk), .RN(rst_n), .Q(
        x_matrix[273]) );
  DFFRHQX1 x_matrix_reg_6__6__1_ ( .D(n4314), .CK(clk), .RN(rst_n), .Q(
        x_matrix[97]) );
  DFFRHQX1 x_matrix_reg_0__2__0_ ( .D(n3483), .CK(clk), .RN(rst_n), .Q(
        x_matrix[720]) );
  DFFRHQX1 x_matrix_reg_2__2__0_ ( .D(n3739), .CK(clk), .RN(rst_n), .Q(
        x_matrix[496]) );
  DFFRHQX1 x_matrix_reg_4__6__0_ ( .D(n4059), .CK(clk), .RN(rst_n), .Q(
        x_matrix[272]) );
  DFFRHQX1 x_matrix_reg_6__6__0_ ( .D(n4315), .CK(clk), .RN(rst_n), .Q(
        x_matrix[96]) );
  DFFRHQX1 x_matrix_reg_0__3__15_ ( .D(n3484), .CK(clk), .RN(rst_n), .Q(
        x_matrix[719]) );
  DFFRHQX1 x_matrix_reg_2__3__15_ ( .D(n3740), .CK(clk), .RN(rst_n), .Q(
        x_matrix[495]) );
  DFFRHQX1 x_matrix_reg_4__7__15_ ( .D(n4060), .CK(clk), .RN(rst_n), .Q(
        x_matrix[271]) );
  DFFRHQX1 x_matrix_reg_6__7__15_ ( .D(n4316), .CK(clk), .RN(rst_n), .Q(
        x_matrix[95]) );
  DFFRHQX1 x_matrix_reg_0__3__14_ ( .D(n3485), .CK(clk), .RN(rst_n), .Q(
        x_matrix[718]) );
  DFFRHQX1 x_matrix_reg_2__3__14_ ( .D(n3741), .CK(clk), .RN(rst_n), .Q(
        x_matrix[494]) );
  DFFRHQX1 x_matrix_reg_4__7__14_ ( .D(n4061), .CK(clk), .RN(rst_n), .Q(
        x_matrix[270]) );
  DFFRHQX1 x_matrix_reg_6__7__14_ ( .D(n4317), .CK(clk), .RN(rst_n), .Q(
        x_matrix[94]) );
  DFFRHQX1 x_matrix_reg_0__3__13_ ( .D(n3486), .CK(clk), .RN(rst_n), .Q(
        x_matrix[717]) );
  DFFRHQX1 x_matrix_reg_2__3__13_ ( .D(n3742), .CK(clk), .RN(rst_n), .Q(
        x_matrix[493]) );
  DFFRHQX1 x_matrix_reg_4__7__13_ ( .D(n4062), .CK(clk), .RN(rst_n), .Q(
        x_matrix[269]) );
  DFFRHQX1 x_matrix_reg_6__7__13_ ( .D(n4318), .CK(clk), .RN(rst_n), .Q(
        x_matrix[93]) );
  DFFRHQX1 x_matrix_reg_0__3__12_ ( .D(n3487), .CK(clk), .RN(rst_n), .Q(
        x_matrix[716]) );
  DFFRHQX1 x_matrix_reg_2__3__12_ ( .D(n3743), .CK(clk), .RN(rst_n), .Q(
        x_matrix[492]) );
  DFFRHQX1 x_matrix_reg_4__7__12_ ( .D(n4063), .CK(clk), .RN(rst_n), .Q(
        x_matrix[268]) );
  DFFRHQX1 x_matrix_reg_6__7__12_ ( .D(n4319), .CK(clk), .RN(rst_n), .Q(
        x_matrix[92]) );
  DFFRHQX1 x_matrix_reg_0__3__11_ ( .D(n3488), .CK(clk), .RN(rst_n), .Q(
        x_matrix[715]) );
  DFFRHQX1 x_matrix_reg_2__3__11_ ( .D(n3744), .CK(clk), .RN(rst_n), .Q(
        x_matrix[491]) );
  DFFRHQX1 x_matrix_reg_4__7__11_ ( .D(n4064), .CK(clk), .RN(rst_n), .Q(
        x_matrix[267]) );
  DFFRHQX1 x_matrix_reg_6__7__11_ ( .D(n4320), .CK(clk), .RN(rst_n), .Q(
        x_matrix[91]) );
  DFFRHQX1 x_matrix_reg_0__3__10_ ( .D(n3489), .CK(clk), .RN(rst_n), .Q(
        x_matrix[714]) );
  DFFRHQX1 x_matrix_reg_2__3__10_ ( .D(n3745), .CK(clk), .RN(rst_n), .Q(
        x_matrix[490]) );
  DFFRHQX1 x_matrix_reg_4__7__10_ ( .D(n4065), .CK(clk), .RN(rst_n), .Q(
        x_matrix[266]) );
  DFFRHQX1 x_matrix_reg_6__7__10_ ( .D(n4321), .CK(clk), .RN(rst_n), .Q(
        x_matrix[90]) );
  DFFRHQX1 x_matrix_reg_0__3__0_ ( .D(n3499), .CK(clk), .RN(rst_n), .Q(
        x_matrix[704]) );
  DFFRHQX1 x_matrix_reg_2__3__0_ ( .D(n3755), .CK(clk), .RN(rst_n), .Q(
        x_matrix[480]) );
  DFFRHQX1 x_matrix_reg_4__7__0_ ( .D(n4075), .CK(clk), .RN(rst_n), .Q(
        x_matrix[256]) );
  DFFRHQX1 x_matrix_reg_6__7__0_ ( .D(n4331), .CK(clk), .RN(rst_n), .Q(
        x_matrix[80]) );
  DFFRHQX1 x_matrix_reg_1__3__9_ ( .D(n3618), .CK(clk), .RN(rst_n), .Q(
        x_matrix[601]) );
  DFFRHQX1 x_matrix_reg_3__3__9_ ( .D(n3874), .CK(clk), .RN(rst_n), .Q(
        x_matrix[393]) );
  DFFRHQX1 x_matrix_reg_5__7__9_ ( .D(n4194), .CK(clk), .RN(rst_n), .Q(
        x_matrix[169]) );
  DFFRHQX1 x_matrix_reg_7__7__9_ ( .D(n4450), .CK(clk), .RN(rst_n), .Q(
        x_matrix[9]) );
  DFFRHQX1 x_matrix_reg_1__3__8_ ( .D(n3619), .CK(clk), .RN(rst_n), .Q(
        x_matrix[600]) );
  DFFRHQX1 x_matrix_reg_3__3__8_ ( .D(n3875), .CK(clk), .RN(rst_n), .Q(
        x_matrix[392]) );
  DFFRHQX1 x_matrix_reg_5__7__8_ ( .D(n4195), .CK(clk), .RN(rst_n), .Q(
        x_matrix[168]) );
  DFFRHQX1 x_matrix_reg_7__7__8_ ( .D(n4451), .CK(clk), .RN(rst_n), .Q(
        x_matrix[8]) );
  DFFRHQX1 x_matrix_reg_1__3__7_ ( .D(n3620), .CK(clk), .RN(rst_n), .Q(
        x_matrix[599]) );
  DFFRHQX1 x_matrix_reg_3__3__7_ ( .D(n3876), .CK(clk), .RN(rst_n), .Q(
        x_matrix[391]) );
  DFFRHQX1 x_matrix_reg_5__7__7_ ( .D(n4196), .CK(clk), .RN(rst_n), .Q(
        x_matrix[167]) );
  DFFRHQX1 x_matrix_reg_7__7__7_ ( .D(n4452), .CK(clk), .RN(rst_n), .Q(
        x_matrix[7]) );
  DFFRHQX1 x_matrix_reg_1__3__6_ ( .D(n3621), .CK(clk), .RN(rst_n), .Q(
        x_matrix[598]) );
  DFFRHQX1 x_matrix_reg_3__3__6_ ( .D(n3877), .CK(clk), .RN(rst_n), .Q(
        x_matrix[390]) );
  DFFRHQX1 x_matrix_reg_5__7__6_ ( .D(n4197), .CK(clk), .RN(rst_n), .Q(
        x_matrix[166]) );
  DFFRHQX1 x_matrix_reg_7__7__6_ ( .D(n4453), .CK(clk), .RN(rst_n), .Q(
        x_matrix[6]) );
  DFFRHQX1 x_matrix_reg_1__4__15_ ( .D(n3628), .CK(clk), .RN(rst_n), .Q(
        x_matrix[591]) );
  DFFRHQX1 x_matrix_reg_3__0__15_ ( .D(n3820), .CK(clk), .RN(rst_n), .Q(
        x_matrix[447]) );
  DFFRHQX1 x_matrix_reg_3__4__15_ ( .D(n3884), .CK(clk), .RN(rst_n), .Q(
        x_matrix[383]) );
  DFFRHQX1 x_matrix_reg_1__4__14_ ( .D(n3629), .CK(clk), .RN(rst_n), .Q(
        x_matrix[590]) );
  DFFRHQX1 x_matrix_reg_3__0__14_ ( .D(n3821), .CK(clk), .RN(rst_n), .Q(
        x_matrix[446]) );
  DFFRHQX1 x_matrix_reg_3__4__14_ ( .D(n3885), .CK(clk), .RN(rst_n), .Q(
        x_matrix[382]) );
  DFFRHQX1 x_matrix_reg_1__4__13_ ( .D(n3630), .CK(clk), .RN(rst_n), .Q(
        x_matrix[589]) );
  DFFRHQX1 x_matrix_reg_3__0__13_ ( .D(n3822), .CK(clk), .RN(rst_n), .Q(
        x_matrix[445]) );
  DFFRHQX1 x_matrix_reg_3__4__13_ ( .D(n3886), .CK(clk), .RN(rst_n), .Q(
        x_matrix[381]) );
  DFFRHQX1 x_matrix_reg_1__4__12_ ( .D(n3631), .CK(clk), .RN(rst_n), .Q(
        x_matrix[588]) );
  DFFRHQX1 x_matrix_reg_3__0__12_ ( .D(n3823), .CK(clk), .RN(rst_n), .Q(
        x_matrix[444]) );
  DFFRHQX1 x_matrix_reg_3__4__12_ ( .D(n3887), .CK(clk), .RN(rst_n), .Q(
        x_matrix[380]) );
  DFFRHQX1 x_matrix_reg_1__3__5_ ( .D(n3622), .CK(clk), .RN(rst_n), .Q(
        x_matrix[597]) );
  DFFRHQX1 x_matrix_reg_3__3__5_ ( .D(n3878), .CK(clk), .RN(rst_n), .Q(
        x_matrix[389]) );
  DFFRHQX1 x_matrix_reg_5__7__5_ ( .D(n4198), .CK(clk), .RN(rst_n), .Q(
        x_matrix[165]) );
  DFFRHQX1 x_matrix_reg_7__7__5_ ( .D(n4454), .CK(clk), .RN(rst_n), .Q(
        x_matrix[5]) );
  DFFRHQX1 x_matrix_reg_1__4__11_ ( .D(n3632), .CK(clk), .RN(rst_n), .Q(
        x_matrix[587]) );
  DFFRHQX1 x_matrix_reg_3__0__11_ ( .D(n3824), .CK(clk), .RN(rst_n), .Q(
        x_matrix[443]) );
  DFFRHQX1 x_matrix_reg_3__4__11_ ( .D(n3888), .CK(clk), .RN(rst_n), .Q(
        x_matrix[379]) );
  DFFRHQX1 x_matrix_reg_1__4__10_ ( .D(n3633), .CK(clk), .RN(rst_n), .Q(
        x_matrix[586]) );
  DFFRHQX1 x_matrix_reg_3__0__10_ ( .D(n3825), .CK(clk), .RN(rst_n), .Q(
        x_matrix[442]) );
  DFFRHQX1 x_matrix_reg_3__4__10_ ( .D(n3889), .CK(clk), .RN(rst_n), .Q(
        x_matrix[378]) );
  DFFRHQX1 x_matrix_reg_1__4__9_ ( .D(n3634), .CK(clk), .RN(rst_n), .Q(
        x_matrix[585]) );
  DFFRHQX1 x_matrix_reg_3__0__9_ ( .D(n3826), .CK(clk), .RN(rst_n), .Q(
        x_matrix[441]) );
  DFFRHQX1 x_matrix_reg_3__4__9_ ( .D(n3890), .CK(clk), .RN(rst_n), .Q(
        x_matrix[377]) );
  DFFRHQX1 x_matrix_reg_1__4__8_ ( .D(n3635), .CK(clk), .RN(rst_n), .Q(
        x_matrix[584]) );
  DFFRHQX1 x_matrix_reg_3__0__8_ ( .D(n3827), .CK(clk), .RN(rst_n), .Q(
        x_matrix[440]) );
  DFFRHQX1 x_matrix_reg_3__4__8_ ( .D(n3891), .CK(clk), .RN(rst_n), .Q(
        x_matrix[376]) );
  DFFRHQX1 x_matrix_reg_1__4__7_ ( .D(n3636), .CK(clk), .RN(rst_n), .Q(
        x_matrix[583]) );
  DFFRHQX1 x_matrix_reg_3__0__7_ ( .D(n3828), .CK(clk), .RN(rst_n), .Q(
        x_matrix[439]) );
  DFFRHQX1 x_matrix_reg_3__4__7_ ( .D(n3892), .CK(clk), .RN(rst_n), .Q(
        x_matrix[375]) );
  DFFRHQX1 x_matrix_reg_1__4__6_ ( .D(n3637), .CK(clk), .RN(rst_n), .Q(
        x_matrix[582]) );
  DFFRHQX1 x_matrix_reg_3__0__6_ ( .D(n3829), .CK(clk), .RN(rst_n), .Q(
        x_matrix[438]) );
  DFFRHQX1 x_matrix_reg_3__4__6_ ( .D(n3893), .CK(clk), .RN(rst_n), .Q(
        x_matrix[374]) );
  DFFRHQX1 x_matrix_reg_1__4__5_ ( .D(n3638), .CK(clk), .RN(rst_n), .Q(
        x_matrix[581]) );
  DFFRHQX1 x_matrix_reg_3__0__5_ ( .D(n3830), .CK(clk), .RN(rst_n), .Q(
        x_matrix[437]) );
  DFFRHQX1 x_matrix_reg_3__4__5_ ( .D(n3894), .CK(clk), .RN(rst_n), .Q(
        x_matrix[373]) );
  DFFRHQX1 x_matrix_reg_1__4__4_ ( .D(n3639), .CK(clk), .RN(rst_n), .Q(
        x_matrix[580]) );
  DFFRHQX1 x_matrix_reg_3__0__4_ ( .D(n3831), .CK(clk), .RN(rst_n), .Q(
        x_matrix[436]) );
  DFFRHQX1 x_matrix_reg_3__4__4_ ( .D(n3895), .CK(clk), .RN(rst_n), .Q(
        x_matrix[372]) );
  DFFRHQX1 x_matrix_reg_1__4__3_ ( .D(n3640), .CK(clk), .RN(rst_n), .Q(
        x_matrix[579]) );
  DFFRHQX1 x_matrix_reg_3__0__3_ ( .D(n3832), .CK(clk), .RN(rst_n), .Q(
        x_matrix[435]) );
  DFFRHQX1 x_matrix_reg_3__4__3_ ( .D(n3896), .CK(clk), .RN(rst_n), .Q(
        x_matrix[371]) );
  DFFRHQX1 x_matrix_reg_1__4__2_ ( .D(n3641), .CK(clk), .RN(rst_n), .Q(
        x_matrix[578]) );
  DFFRHQX1 x_matrix_reg_3__0__2_ ( .D(n3833), .CK(clk), .RN(rst_n), .Q(
        x_matrix[434]) );
  DFFRHQX1 x_matrix_reg_3__4__2_ ( .D(n3897), .CK(clk), .RN(rst_n), .Q(
        x_matrix[370]) );
  DFFRHQX1 x_matrix_reg_1__3__4_ ( .D(n3623), .CK(clk), .RN(rst_n), .Q(
        x_matrix[596]) );
  DFFRHQX1 x_matrix_reg_3__3__4_ ( .D(n3879), .CK(clk), .RN(rst_n), .Q(
        x_matrix[388]) );
  DFFRHQX1 x_matrix_reg_5__7__4_ ( .D(n4199), .CK(clk), .RN(rst_n), .Q(
        x_matrix[164]) );
  DFFRHQX1 x_matrix_reg_7__7__4_ ( .D(n4455), .CK(clk), .RN(rst_n), .Q(
        x_matrix[4]) );
  DFFRHQX1 x_matrix_reg_1__4__1_ ( .D(n3642), .CK(clk), .RN(rst_n), .Q(
        x_matrix[577]) );
  DFFRHQX1 x_matrix_reg_3__0__1_ ( .D(n3834), .CK(clk), .RN(rst_n), .Q(
        x_matrix[433]) );
  DFFRHQX1 x_matrix_reg_3__4__1_ ( .D(n3898), .CK(clk), .RN(rst_n), .Q(
        x_matrix[369]) );
  DFFRHQX1 x_matrix_reg_1__4__0_ ( .D(n3643), .CK(clk), .RN(rst_n), .Q(
        x_matrix[576]) );
  DFFRHQX1 x_matrix_reg_3__0__0_ ( .D(n3835), .CK(clk), .RN(rst_n), .Q(
        x_matrix[432]) );
  DFFRHQX1 x_matrix_reg_3__4__0_ ( .D(n3899), .CK(clk), .RN(rst_n), .Q(
        x_matrix[368]) );
  DFFRHQX1 x_matrix_reg_3__1__15_ ( .D(n3836), .CK(clk), .RN(rst_n), .Q(
        x_matrix[431]) );
  DFFRHQX1 x_matrix_reg_5__5__15_ ( .D(n4156), .CK(clk), .RN(rst_n), .Q(
        x_matrix[207]) );
  DFFRHQX1 x_matrix_reg_7__5__15_ ( .D(n4412), .CK(clk), .RN(rst_n), .Q(
        x_matrix[47]) );
  DFFRHQX1 x_matrix_reg_3__1__14_ ( .D(n3837), .CK(clk), .RN(rst_n), .Q(
        x_matrix[430]) );
  DFFRHQX1 x_matrix_reg_5__5__14_ ( .D(n4157), .CK(clk), .RN(rst_n), .Q(
        x_matrix[206]) );
  DFFRHQX1 x_matrix_reg_7__5__14_ ( .D(n4413), .CK(clk), .RN(rst_n), .Q(
        x_matrix[46]) );
  DFFRHQX1 x_matrix_reg_3__1__13_ ( .D(n3838), .CK(clk), .RN(rst_n), .Q(
        x_matrix[429]) );
  DFFRHQX1 x_matrix_reg_5__5__13_ ( .D(n4158), .CK(clk), .RN(rst_n), .Q(
        x_matrix[205]) );
  DFFRHQX1 x_matrix_reg_7__5__13_ ( .D(n4414), .CK(clk), .RN(rst_n), .Q(
        x_matrix[45]) );
  DFFRHQX1 x_matrix_reg_3__1__12_ ( .D(n3839), .CK(clk), .RN(rst_n), .Q(
        x_matrix[428]) );
  DFFRHQX1 x_matrix_reg_5__5__12_ ( .D(n4159), .CK(clk), .RN(rst_n), .Q(
        x_matrix[204]) );
  DFFRHQX1 x_matrix_reg_7__5__12_ ( .D(n4415), .CK(clk), .RN(rst_n), .Q(
        x_matrix[44]) );
  DFFRHQX1 x_matrix_reg_3__1__11_ ( .D(n3840), .CK(clk), .RN(rst_n), .Q(
        x_matrix[427]) );
  DFFRHQX1 x_matrix_reg_5__5__11_ ( .D(n4160), .CK(clk), .RN(rst_n), .Q(
        x_matrix[203]) );
  DFFRHQX1 x_matrix_reg_7__5__11_ ( .D(n4416), .CK(clk), .RN(rst_n), .Q(
        x_matrix[43]) );
  DFFRHQX1 x_matrix_reg_3__1__10_ ( .D(n3841), .CK(clk), .RN(rst_n), .Q(
        x_matrix[426]) );
  DFFRHQX1 x_matrix_reg_5__5__10_ ( .D(n4161), .CK(clk), .RN(rst_n), .Q(
        x_matrix[202]) );
  DFFRHQX1 x_matrix_reg_7__5__10_ ( .D(n4417), .CK(clk), .RN(rst_n), .Q(
        x_matrix[42]) );
  DFFRHQX1 x_matrix_reg_3__1__9_ ( .D(n3842), .CK(clk), .RN(rst_n), .Q(
        x_matrix[425]) );
  DFFRHQX1 x_matrix_reg_5__5__9_ ( .D(n4162), .CK(clk), .RN(rst_n), .Q(
        x_matrix[201]) );
  DFFRHQX1 x_matrix_reg_7__5__9_ ( .D(n4418), .CK(clk), .RN(rst_n), .Q(
        x_matrix[41]) );
  DFFRHQX1 x_matrix_reg_3__1__8_ ( .D(n3843), .CK(clk), .RN(rst_n), .Q(
        x_matrix[424]) );
  DFFRHQX1 x_matrix_reg_5__5__8_ ( .D(n4163), .CK(clk), .RN(rst_n), .Q(
        x_matrix[200]) );
  DFFRHQX1 x_matrix_reg_7__5__8_ ( .D(n4419), .CK(clk), .RN(rst_n), .Q(
        x_matrix[40]) );
  DFFRHQX1 x_matrix_reg_1__3__3_ ( .D(n3624), .CK(clk), .RN(rst_n), .Q(
        x_matrix[595]) );
  DFFRHQX1 x_matrix_reg_3__3__3_ ( .D(n3880), .CK(clk), .RN(rst_n), .Q(
        x_matrix[387]) );
  DFFRHQX1 x_matrix_reg_5__7__3_ ( .D(n4200), .CK(clk), .RN(rst_n), .Q(
        x_matrix[163]) );
  DFFRHQX1 x_matrix_reg_7__7__3_ ( .D(n4456), .CK(clk), .RN(rst_n), .Q(
        x_matrix[3]) );
  DFFRHQX1 x_matrix_reg_3__1__7_ ( .D(n3844), .CK(clk), .RN(rst_n), .Q(
        x_matrix[423]) );
  DFFRHQX1 x_matrix_reg_5__5__7_ ( .D(n4164), .CK(clk), .RN(rst_n), .Q(
        x_matrix[199]) );
  DFFRHQX1 x_matrix_reg_7__5__7_ ( .D(n4420), .CK(clk), .RN(rst_n), .Q(
        x_matrix[39]) );
  DFFRHQX1 x_matrix_reg_3__1__6_ ( .D(n3845), .CK(clk), .RN(rst_n), .Q(
        x_matrix[422]) );
  DFFRHQX1 x_matrix_reg_5__5__6_ ( .D(n4165), .CK(clk), .RN(rst_n), .Q(
        x_matrix[198]) );
  DFFRHQX1 x_matrix_reg_7__5__6_ ( .D(n4421), .CK(clk), .RN(rst_n), .Q(
        x_matrix[38]) );
  DFFRHQX1 x_matrix_reg_3__1__5_ ( .D(n3846), .CK(clk), .RN(rst_n), .Q(
        x_matrix[421]) );
  DFFRHQX1 x_matrix_reg_5__5__5_ ( .D(n4166), .CK(clk), .RN(rst_n), .Q(
        x_matrix[197]) );
  DFFRHQX1 x_matrix_reg_7__5__5_ ( .D(n4422), .CK(clk), .RN(rst_n), .Q(
        x_matrix[37]) );
  DFFRHQX1 x_matrix_reg_3__1__4_ ( .D(n3847), .CK(clk), .RN(rst_n), .Q(
        x_matrix[420]) );
  DFFRHQX1 x_matrix_reg_5__5__4_ ( .D(n4167), .CK(clk), .RN(rst_n), .Q(
        x_matrix[196]) );
  DFFRHQX1 x_matrix_reg_7__5__4_ ( .D(n4423), .CK(clk), .RN(rst_n), .Q(
        x_matrix[36]) );
  DFFRHQX1 x_matrix_reg_3__1__3_ ( .D(n3848), .CK(clk), .RN(rst_n), .Q(
        x_matrix[419]) );
  DFFRHQX1 x_matrix_reg_5__5__3_ ( .D(n4168), .CK(clk), .RN(rst_n), .Q(
        x_matrix[195]) );
  DFFRHQX1 x_matrix_reg_7__5__3_ ( .D(n4424), .CK(clk), .RN(rst_n), .Q(
        x_matrix[35]) );
  DFFRHQX1 x_matrix_reg_3__1__2_ ( .D(n3849), .CK(clk), .RN(rst_n), .Q(
        x_matrix[418]) );
  DFFRHQX1 x_matrix_reg_5__5__2_ ( .D(n4169), .CK(clk), .RN(rst_n), .Q(
        x_matrix[194]) );
  DFFRHQX1 x_matrix_reg_7__5__2_ ( .D(n4425), .CK(clk), .RN(rst_n), .Q(
        x_matrix[34]) );
  DFFRHQX1 x_matrix_reg_3__1__1_ ( .D(n3850), .CK(clk), .RN(rst_n), .Q(
        x_matrix[417]) );
  DFFRHQX1 x_matrix_reg_5__5__1_ ( .D(n4170), .CK(clk), .RN(rst_n), .Q(
        x_matrix[193]) );
  DFFRHQX1 x_matrix_reg_7__5__1_ ( .D(n4426), .CK(clk), .RN(rst_n), .Q(
        x_matrix[33]) );
  DFFRHQX1 x_matrix_reg_3__1__0_ ( .D(n3851), .CK(clk), .RN(rst_n), .Q(
        x_matrix[416]) );
  DFFRHQX1 x_matrix_reg_5__5__0_ ( .D(n4171), .CK(clk), .RN(rst_n), .Q(
        x_matrix[192]) );
  DFFRHQX1 x_matrix_reg_7__5__0_ ( .D(n4427), .CK(clk), .RN(rst_n), .Q(
        x_matrix[32]) );
  DFFRHQX1 x_matrix_reg_1__2__15_ ( .D(n3596), .CK(clk), .RN(rst_n), .Q(
        x_matrix[623]) );
  DFFRHQX1 x_matrix_reg_3__2__15_ ( .D(n3852), .CK(clk), .RN(rst_n), .Q(
        x_matrix[415]) );
  DFFRHQX1 x_matrix_reg_5__6__15_ ( .D(n4172), .CK(clk), .RN(rst_n), .Q(
        x_matrix[191]) );
  DFFRHQX1 x_matrix_reg_7__6__15_ ( .D(n4428), .CK(clk), .RN(rst_n), .Q(
        x_matrix[31]) );
  DFFRHQX1 x_matrix_reg_1__2__14_ ( .D(n3597), .CK(clk), .RN(rst_n), .Q(
        x_matrix[622]) );
  DFFRHQX1 x_matrix_reg_3__2__14_ ( .D(n3853), .CK(clk), .RN(rst_n), .Q(
        x_matrix[414]) );
  DFFRHQX1 x_matrix_reg_5__6__14_ ( .D(n4173), .CK(clk), .RN(rst_n), .Q(
        x_matrix[190]) );
  DFFRHQX1 x_matrix_reg_7__6__14_ ( .D(n4429), .CK(clk), .RN(rst_n), .Q(
        x_matrix[30]) );
  DFFRHQX1 x_matrix_reg_1__3__2_ ( .D(n3625), .CK(clk), .RN(rst_n), .Q(
        x_matrix[594]) );
  DFFRHQX1 x_matrix_reg_3__3__2_ ( .D(n3881), .CK(clk), .RN(rst_n), .Q(
        x_matrix[386]) );
  DFFRHQX1 x_matrix_reg_5__7__2_ ( .D(n4201), .CK(clk), .RN(rst_n), .Q(
        x_matrix[162]) );
  DFFRHQX1 x_matrix_reg_7__7__2_ ( .D(n4457), .CK(clk), .RN(rst_n), .Q(
        x_matrix[2]) );
  DFFRHQX1 x_matrix_reg_1__2__13_ ( .D(n3598), .CK(clk), .RN(rst_n), .Q(
        x_matrix[621]) );
  DFFRHQX1 x_matrix_reg_3__2__13_ ( .D(n3854), .CK(clk), .RN(rst_n), .Q(
        x_matrix[413]) );
  DFFRHQX1 x_matrix_reg_5__6__13_ ( .D(n4174), .CK(clk), .RN(rst_n), .Q(
        x_matrix[189]) );
  DFFRHQX1 x_matrix_reg_7__6__13_ ( .D(n4430), .CK(clk), .RN(rst_n), .Q(
        x_matrix[29]) );
  DFFRHQX1 x_matrix_reg_1__2__12_ ( .D(n3599), .CK(clk), .RN(rst_n), .Q(
        x_matrix[620]) );
  DFFRHQX1 x_matrix_reg_3__2__12_ ( .D(n3855), .CK(clk), .RN(rst_n), .Q(
        x_matrix[412]) );
  DFFRHQX1 x_matrix_reg_5__6__12_ ( .D(n4175), .CK(clk), .RN(rst_n), .Q(
        x_matrix[188]) );
  DFFRHQX1 x_matrix_reg_7__6__12_ ( .D(n4431), .CK(clk), .RN(rst_n), .Q(
        x_matrix[28]) );
  DFFRHQX1 x_matrix_reg_1__2__11_ ( .D(n3600), .CK(clk), .RN(rst_n), .Q(
        x_matrix[619]) );
  DFFRHQX1 x_matrix_reg_3__2__11_ ( .D(n3856), .CK(clk), .RN(rst_n), .Q(
        x_matrix[411]) );
  DFFRHQX1 x_matrix_reg_5__6__11_ ( .D(n4176), .CK(clk), .RN(rst_n), .Q(
        x_matrix[187]) );
  DFFRHQX1 x_matrix_reg_7__6__11_ ( .D(n4432), .CK(clk), .RN(rst_n), .Q(
        x_matrix[27]) );
  DFFRHQX1 x_matrix_reg_1__2__10_ ( .D(n3601), .CK(clk), .RN(rst_n), .Q(
        x_matrix[618]) );
  DFFRHQX1 x_matrix_reg_3__2__10_ ( .D(n3857), .CK(clk), .RN(rst_n), .Q(
        x_matrix[410]) );
  DFFRHQX1 x_matrix_reg_5__6__10_ ( .D(n4177), .CK(clk), .RN(rst_n), .Q(
        x_matrix[186]) );
  DFFRHQX1 x_matrix_reg_7__6__10_ ( .D(n4433), .CK(clk), .RN(rst_n), .Q(
        x_matrix[26]) );
  DFFRHQX1 x_matrix_reg_1__2__9_ ( .D(n3602), .CK(clk), .RN(rst_n), .Q(
        x_matrix[617]) );
  DFFRHQX1 x_matrix_reg_3__2__9_ ( .D(n3858), .CK(clk), .RN(rst_n), .Q(
        x_matrix[409]) );
  DFFRHQX1 x_matrix_reg_5__6__9_ ( .D(n4178), .CK(clk), .RN(rst_n), .Q(
        x_matrix[185]) );
  DFFRHQX1 x_matrix_reg_7__6__9_ ( .D(n4434), .CK(clk), .RN(rst_n), .Q(
        x_matrix[25]) );
  DFFRHQX1 x_matrix_reg_1__2__8_ ( .D(n3603), .CK(clk), .RN(rst_n), .Q(
        x_matrix[616]) );
  DFFRHQX1 x_matrix_reg_3__2__8_ ( .D(n3859), .CK(clk), .RN(rst_n), .Q(
        x_matrix[408]) );
  DFFRHQX1 x_matrix_reg_5__6__8_ ( .D(n4179), .CK(clk), .RN(rst_n), .Q(
        x_matrix[184]) );
  DFFRHQX1 x_matrix_reg_7__6__8_ ( .D(n4435), .CK(clk), .RN(rst_n), .Q(
        x_matrix[24]) );
  DFFRHQX1 x_matrix_reg_1__2__7_ ( .D(n3604), .CK(clk), .RN(rst_n), .Q(
        x_matrix[615]) );
  DFFRHQX1 x_matrix_reg_3__2__7_ ( .D(n3860), .CK(clk), .RN(rst_n), .Q(
        x_matrix[407]) );
  DFFRHQX1 x_matrix_reg_5__6__7_ ( .D(n4180), .CK(clk), .RN(rst_n), .Q(
        x_matrix[183]) );
  DFFRHQX1 x_matrix_reg_7__6__7_ ( .D(n4436), .CK(clk), .RN(rst_n), .Q(
        x_matrix[23]) );
  DFFRHQX1 x_matrix_reg_1__2__6_ ( .D(n3605), .CK(clk), .RN(rst_n), .Q(
        x_matrix[614]) );
  DFFRHQX1 x_matrix_reg_3__2__6_ ( .D(n3861), .CK(clk), .RN(rst_n), .Q(
        x_matrix[406]) );
  DFFRHQX1 x_matrix_reg_5__6__6_ ( .D(n4181), .CK(clk), .RN(rst_n), .Q(
        x_matrix[182]) );
  DFFRHQX1 x_matrix_reg_7__6__6_ ( .D(n4437), .CK(clk), .RN(rst_n), .Q(
        x_matrix[22]) );
  DFFRHQX1 x_matrix_reg_1__2__5_ ( .D(n3606), .CK(clk), .RN(rst_n), .Q(
        x_matrix[613]) );
  DFFRHQX1 x_matrix_reg_3__2__5_ ( .D(n3862), .CK(clk), .RN(rst_n), .Q(
        x_matrix[405]) );
  DFFRHQX1 x_matrix_reg_5__6__5_ ( .D(n4182), .CK(clk), .RN(rst_n), .Q(
        x_matrix[181]) );
  DFFRHQX1 x_matrix_reg_7__6__5_ ( .D(n4438), .CK(clk), .RN(rst_n), .Q(
        x_matrix[21]) );
  DFFRHQX1 x_matrix_reg_1__2__4_ ( .D(n3607), .CK(clk), .RN(rst_n), .Q(
        x_matrix[612]) );
  DFFRHQX1 x_matrix_reg_3__2__4_ ( .D(n3863), .CK(clk), .RN(rst_n), .Q(
        x_matrix[404]) );
  DFFRHQX1 x_matrix_reg_5__6__4_ ( .D(n4183), .CK(clk), .RN(rst_n), .Q(
        x_matrix[180]) );
  DFFRHQX1 x_matrix_reg_7__6__4_ ( .D(n4439), .CK(clk), .RN(rst_n), .Q(
        x_matrix[20]) );
  DFFRHQX1 x_matrix_reg_1__3__1_ ( .D(n3626), .CK(clk), .RN(rst_n), .Q(
        x_matrix[593]) );
  DFFRHQX1 x_matrix_reg_3__3__1_ ( .D(n3882), .CK(clk), .RN(rst_n), .Q(
        x_matrix[385]) );
  DFFRHQX1 x_matrix_reg_5__7__1_ ( .D(n4202), .CK(clk), .RN(rst_n), .Q(
        x_matrix[161]) );
  DFFRHQX1 x_matrix_reg_7__7__1_ ( .D(n4458), .CK(clk), .RN(rst_n), .Q(
        x_matrix[1]) );
  DFFRHQX1 x_matrix_reg_1__2__3_ ( .D(n3608), .CK(clk), .RN(rst_n), .Q(
        x_matrix[611]) );
  DFFRHQX1 x_matrix_reg_3__2__3_ ( .D(n3864), .CK(clk), .RN(rst_n), .Q(
        x_matrix[403]) );
  DFFRHQX1 x_matrix_reg_5__6__3_ ( .D(n4184), .CK(clk), .RN(rst_n), .Q(
        x_matrix[179]) );
  DFFRHQX1 x_matrix_reg_7__6__3_ ( .D(n4440), .CK(clk), .RN(rst_n), .Q(
        x_matrix[19]) );
  DFFRHQX1 x_matrix_reg_1__2__2_ ( .D(n3609), .CK(clk), .RN(rst_n), .Q(
        x_matrix[610]) );
  DFFRHQX1 x_matrix_reg_3__2__2_ ( .D(n3865), .CK(clk), .RN(rst_n), .Q(
        x_matrix[402]) );
  DFFRHQX1 x_matrix_reg_5__6__2_ ( .D(n4185), .CK(clk), .RN(rst_n), .Q(
        x_matrix[178]) );
  DFFRHQX1 x_matrix_reg_7__6__2_ ( .D(n4441), .CK(clk), .RN(rst_n), .Q(
        x_matrix[18]) );
  DFFRHQX1 x_matrix_reg_1__2__1_ ( .D(n3610), .CK(clk), .RN(rst_n), .Q(
        x_matrix[609]) );
  DFFRHQX1 x_matrix_reg_3__2__1_ ( .D(n3866), .CK(clk), .RN(rst_n), .Q(
        x_matrix[401]) );
  DFFRHQX1 x_matrix_reg_5__6__1_ ( .D(n4186), .CK(clk), .RN(rst_n), .Q(
        x_matrix[177]) );
  DFFRHQX1 x_matrix_reg_7__6__1_ ( .D(n4442), .CK(clk), .RN(rst_n), .Q(
        x_matrix[17]) );
  DFFRHQX1 x_matrix_reg_1__2__0_ ( .D(n3611), .CK(clk), .RN(rst_n), .Q(
        x_matrix[608]) );
  DFFRHQX1 x_matrix_reg_3__2__0_ ( .D(n3867), .CK(clk), .RN(rst_n), .Q(
        x_matrix[400]) );
  DFFRHQX1 x_matrix_reg_5__6__0_ ( .D(n4187), .CK(clk), .RN(rst_n), .Q(
        x_matrix[176]) );
  DFFRHQX1 x_matrix_reg_7__6__0_ ( .D(n4443), .CK(clk), .RN(rst_n), .Q(
        x_matrix[16]) );
  DFFRHQX1 x_matrix_reg_1__3__15_ ( .D(n3612), .CK(clk), .RN(rst_n), .Q(
        x_matrix[607]) );
  DFFRHQX1 x_matrix_reg_3__3__15_ ( .D(n3868), .CK(clk), .RN(rst_n), .Q(
        x_matrix[399]) );
  DFFRHQX1 x_matrix_reg_5__7__15_ ( .D(n4188), .CK(clk), .RN(rst_n), .Q(
        x_matrix[175]) );
  DFFRHQX1 x_matrix_reg_7__7__15_ ( .D(n4444), .CK(clk), .RN(rst_n), .Q(
        x_matrix[15]) );
  DFFRHQX1 x_matrix_reg_1__3__14_ ( .D(n3613), .CK(clk), .RN(rst_n), .Q(
        x_matrix[606]) );
  DFFRHQX1 x_matrix_reg_3__3__14_ ( .D(n3869), .CK(clk), .RN(rst_n), .Q(
        x_matrix[398]) );
  DFFRHQX1 x_matrix_reg_5__7__14_ ( .D(n4189), .CK(clk), .RN(rst_n), .Q(
        x_matrix[174]) );
  DFFRHQX1 x_matrix_reg_7__7__14_ ( .D(n4445), .CK(clk), .RN(rst_n), .Q(
        x_matrix[14]) );
  DFFRHQX1 x_matrix_reg_1__3__13_ ( .D(n3614), .CK(clk), .RN(rst_n), .Q(
        x_matrix[605]) );
  DFFRHQX1 x_matrix_reg_3__3__13_ ( .D(n3870), .CK(clk), .RN(rst_n), .Q(
        x_matrix[397]) );
  DFFRHQX1 x_matrix_reg_5__7__13_ ( .D(n4190), .CK(clk), .RN(rst_n), .Q(
        x_matrix[173]) );
  DFFRHQX1 x_matrix_reg_7__7__13_ ( .D(n4446), .CK(clk), .RN(rst_n), .Q(
        x_matrix[13]) );
  DFFRHQX1 x_matrix_reg_1__3__12_ ( .D(n3615), .CK(clk), .RN(rst_n), .Q(
        x_matrix[604]) );
  DFFRHQX1 x_matrix_reg_3__3__12_ ( .D(n3871), .CK(clk), .RN(rst_n), .Q(
        x_matrix[396]) );
  DFFRHQX1 x_matrix_reg_5__7__12_ ( .D(n4191), .CK(clk), .RN(rst_n), .Q(
        x_matrix[172]) );
  DFFRHQX1 x_matrix_reg_7__7__12_ ( .D(n4447), .CK(clk), .RN(rst_n), .Q(
        x_matrix[12]) );
  DFFRHQX1 x_matrix_reg_1__3__11_ ( .D(n3616), .CK(clk), .RN(rst_n), .Q(
        x_matrix[603]) );
  DFFRHQX1 x_matrix_reg_3__3__11_ ( .D(n3872), .CK(clk), .RN(rst_n), .Q(
        x_matrix[395]) );
  DFFRHQX1 x_matrix_reg_5__7__11_ ( .D(n4192), .CK(clk), .RN(rst_n), .Q(
        x_matrix[171]) );
  DFFRHQX1 x_matrix_reg_7__7__11_ ( .D(n4448), .CK(clk), .RN(rst_n), .Q(
        x_matrix[11]) );
  DFFRHQX1 x_matrix_reg_1__3__10_ ( .D(n3617), .CK(clk), .RN(rst_n), .Q(
        x_matrix[602]) );
  DFFRHQX1 x_matrix_reg_3__3__10_ ( .D(n3873), .CK(clk), .RN(rst_n), .Q(
        x_matrix[394]) );
  DFFRHQX1 x_matrix_reg_5__7__10_ ( .D(n4193), .CK(clk), .RN(rst_n), .Q(
        x_matrix[170]) );
  DFFRHQX1 x_matrix_reg_7__7__10_ ( .D(n4449), .CK(clk), .RN(rst_n), .Q(
        x_matrix[10]) );
  DFFRHQX1 x_matrix_reg_1__3__0_ ( .D(n3627), .CK(clk), .RN(rst_n), .Q(
        x_matrix[592]) );
  DFFRHQX1 x_matrix_reg_3__3__0_ ( .D(n3883), .CK(clk), .RN(rst_n), .Q(
        x_matrix[384]) );
  DFFRHQX1 x_matrix_reg_5__7__0_ ( .D(n4203), .CK(clk), .RN(rst_n), .Q(
        x_matrix[160]) );
  DFFRHQX1 x_matrix_reg_7__7__0_ ( .D(n4459), .CK(clk), .RN(rst_n), .Q(
        x_matrix[0]) );
  DFFRHQX1 c_plus_reg_2_ ( .D(N12568), .CK(clk), .RN(rst_n), .Q(c_plus[2]) );
  DFFSX1 in_addr_cnt_reg_8_ ( .D(n4461), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[8]) );
  DFFRHQX1 in_weight_flag_reg ( .D(n5798), .CK(clk), .RN(rst_n), .Q(
        in_weight_flag) );
  DFFRHQX1 in_matrix_cnt_reg_4_ ( .D(n5796), .CK(clk), .RN(rst_n), .Q(N1276)
         );
  DFFRHQX1 x_matrix_reg_1__1__9_ ( .D(n3586), .CK(clk), .RN(rst_n), .Q(
        x_matrix[633]) );
  DFFRHQX1 x_matrix_reg_1__1__8_ ( .D(n3587), .CK(clk), .RN(rst_n), .Q(
        x_matrix[632]) );
  DFFRHQX1 x_matrix_reg_1__1__7_ ( .D(n3588), .CK(clk), .RN(rst_n), .Q(
        x_matrix[631]) );
  DFFRHQX1 x_matrix_reg_1__1__6_ ( .D(n3589), .CK(clk), .RN(rst_n), .Q(
        x_matrix[630]) );
  DFFRHQX1 x_matrix_reg_1__1__5_ ( .D(n3590), .CK(clk), .RN(rst_n), .Q(
        x_matrix[629]) );
  DFFRHQX1 x_matrix_reg_1__1__4_ ( .D(n3591), .CK(clk), .RN(rst_n), .Q(
        x_matrix[628]) );
  DFFRHQX1 x_matrix_reg_1__1__3_ ( .D(n3592), .CK(clk), .RN(rst_n), .Q(
        x_matrix[627]) );
  DFFRHQX1 x_matrix_reg_1__0__15_ ( .D(n3564), .CK(clk), .RN(rst_n), .Q(
        x_matrix[655]) );
  DFFRHQX1 x_matrix_reg_1__0__14_ ( .D(n3565), .CK(clk), .RN(rst_n), .Q(
        x_matrix[654]) );
  DFFRHQX1 x_matrix_reg_1__1__2_ ( .D(n3593), .CK(clk), .RN(rst_n), .Q(
        x_matrix[626]) );
  DFFRHQX1 x_matrix_reg_1__0__13_ ( .D(n3566), .CK(clk), .RN(rst_n), .Q(
        x_matrix[653]) );
  DFFRHQX1 x_matrix_reg_1__0__12_ ( .D(n3567), .CK(clk), .RN(rst_n), .Q(
        x_matrix[652]) );
  DFFRHQX1 x_matrix_reg_1__0__11_ ( .D(n3568), .CK(clk), .RN(rst_n), .Q(
        x_matrix[651]) );
  DFFRHQX1 x_matrix_reg_1__0__10_ ( .D(n3569), .CK(clk), .RN(rst_n), .Q(
        x_matrix[650]) );
  DFFRHQX1 x_matrix_reg_1__0__9_ ( .D(n3570), .CK(clk), .RN(rst_n), .Q(
        x_matrix[649]) );
  DFFRHQX1 x_matrix_reg_1__0__8_ ( .D(n3571), .CK(clk), .RN(rst_n), .Q(
        x_matrix[648]) );
  DFFRHQX1 x_matrix_reg_1__0__7_ ( .D(n3572), .CK(clk), .RN(rst_n), .Q(
        x_matrix[647]) );
  DFFRHQX1 x_matrix_reg_1__0__6_ ( .D(n3573), .CK(clk), .RN(rst_n), .Q(
        x_matrix[646]) );
  DFFRHQX1 x_matrix_reg_1__0__5_ ( .D(n3574), .CK(clk), .RN(rst_n), .Q(
        x_matrix[645]) );
  DFFRHQX1 x_matrix_reg_1__0__4_ ( .D(n3575), .CK(clk), .RN(rst_n), .Q(
        x_matrix[644]) );
  DFFRHQX1 x_matrix_reg_1__1__1_ ( .D(n3594), .CK(clk), .RN(rst_n), .Q(
        x_matrix[625]) );
  DFFRHQX1 x_matrix_reg_1__0__3_ ( .D(n3576), .CK(clk), .RN(rst_n), .Q(
        x_matrix[643]) );
  DFFRHQX1 x_matrix_reg_1__0__2_ ( .D(n3577), .CK(clk), .RN(rst_n), .Q(
        x_matrix[642]) );
  DFFRHQX1 x_matrix_reg_1__0__1_ ( .D(n3578), .CK(clk), .RN(rst_n), .Q(
        x_matrix[641]) );
  DFFRHQX1 x_matrix_reg_1__0__0_ ( .D(n3579), .CK(clk), .RN(rst_n), .Q(
        x_matrix[640]) );
  DFFRHQX1 x_matrix_reg_1__1__15_ ( .D(n3580), .CK(clk), .RN(rst_n), .Q(
        x_matrix[639]) );
  DFFRHQX1 x_matrix_reg_1__1__14_ ( .D(n3581), .CK(clk), .RN(rst_n), .Q(
        x_matrix[638]) );
  DFFRHQX1 x_matrix_reg_1__1__13_ ( .D(n3582), .CK(clk), .RN(rst_n), .Q(
        x_matrix[637]) );
  DFFRHQX1 x_matrix_reg_1__1__12_ ( .D(n3583), .CK(clk), .RN(rst_n), .Q(
        x_matrix[636]) );
  DFFRHQX1 x_matrix_reg_1__1__11_ ( .D(n3584), .CK(clk), .RN(rst_n), .Q(
        x_matrix[635]) );
  DFFRHQX1 x_matrix_reg_1__1__10_ ( .D(n3585), .CK(clk), .RN(rst_n), .Q(
        x_matrix[634]) );
  DFFRHQX1 x_matrix_reg_1__1__0_ ( .D(n3595), .CK(clk), .RN(rst_n), .Q(
        x_matrix[624]) );
  DFFRHQX1 calweight_addr_reg_8_ ( .D(n5820), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[8]) );
  DFFRHQX1 calin_addr_reg_8_ ( .D(n5811), .CK(clk), .RN(rst_n), .Q(
        calin_addr[8]) );
  DFFRHQX1 c_plus_reg_1_ ( .D(N12567), .CK(clk), .RN(rst_n), .Q(c_plus[1]) );
  DFFRHQX1 c_plus_reg_0_ ( .D(N12566), .CK(clk), .RN(rst_n), .Q(c_plus[0]) );
  DFFRHQX1 cal_out_reg_1__0_ ( .D(n1891), .CK(clk), .RN(rst_n), .Q(
        cal_out[520]) );
  DFFRHQX1 cal_out_reg_3__0_ ( .D(n1971), .CK(clk), .RN(rst_n), .Q(
        cal_out[440]) );
  DFFRHQX1 cal_out_reg_5__0_ ( .D(n2051), .CK(clk), .RN(rst_n), .Q(
        cal_out[360]) );
  DFFRHQX1 cal_out_reg_7__0_ ( .D(n2131), .CK(clk), .RN(rst_n), .Q(
        cal_out[280]) );
  DFFRHQX1 cal_out_reg_11__0_ ( .D(n2291), .CK(clk), .RN(rst_n), .Q(
        cal_out[120]) );
  DFFRHQX1 cal_out_reg_13__0_ ( .D(n2371), .CK(clk), .RN(rst_n), .Q(
        cal_out[40]) );
  DFFRHQX1 cal_out_reg_5__1_ ( .D(n2050), .CK(clk), .RN(rst_n), .Q(
        cal_out[361]) );
  DFFRHQX1 cal_out_reg_11__1_ ( .D(n2290), .CK(clk), .RN(rst_n), .Q(
        cal_out[121]) );
  DFFRHQX1 cal_out_reg_5__3_ ( .D(n2048), .CK(clk), .RN(rst_n), .Q(
        cal_out[363]) );
  DFFRHQX1 cal_out_reg_11__3_ ( .D(n2288), .CK(clk), .RN(rst_n), .Q(
        cal_out[123]) );
  DFFRHQX1 cal_out_reg_1__4_ ( .D(n1887), .CK(clk), .RN(rst_n), .Q(
        cal_out[524]) );
  DFFRHQX1 cal_out_reg_3__4_ ( .D(n1967), .CK(clk), .RN(rst_n), .Q(
        cal_out[444]) );
  DFFRHQX1 cal_out_reg_5__4_ ( .D(n2047), .CK(clk), .RN(rst_n), .Q(
        cal_out[364]) );
  DFFRHQX1 cal_out_reg_7__4_ ( .D(n2127), .CK(clk), .RN(rst_n), .Q(
        cal_out[284]) );
  DFFRHQX1 cal_out_reg_11__4_ ( .D(n2287), .CK(clk), .RN(rst_n), .Q(
        cal_out[124]) );
  DFFRHQX1 cal_out_reg_13__4_ ( .D(n2367), .CK(clk), .RN(rst_n), .Q(
        cal_out[44]) );
  DFFRHQX1 cal_out_reg_5__5_ ( .D(n2046), .CK(clk), .RN(rst_n), .Q(
        cal_out[365]) );
  DFFRHQX1 cal_out_reg_11__5_ ( .D(n2286), .CK(clk), .RN(rst_n), .Q(
        cal_out[125]) );
  DFFRHQX1 cal_out_reg_1__6_ ( .D(n1885), .CK(clk), .RN(rst_n), .Q(
        cal_out[526]) );
  DFFRHQX1 cal_out_reg_3__6_ ( .D(n1965), .CK(clk), .RN(rst_n), .Q(
        cal_out[446]) );
  DFFRHQX1 cal_out_reg_5__6_ ( .D(n2045), .CK(clk), .RN(rst_n), .Q(
        cal_out[366]) );
  DFFRHQX1 cal_out_reg_7__6_ ( .D(n2125), .CK(clk), .RN(rst_n), .Q(
        cal_out[286]) );
  DFFRHQX1 cal_out_reg_11__6_ ( .D(n2285), .CK(clk), .RN(rst_n), .Q(
        cal_out[126]) );
  DFFRHQX1 cal_out_reg_13__6_ ( .D(n2365), .CK(clk), .RN(rst_n), .Q(
        cal_out[46]) );
  DFFRHQX1 cal_out_reg_5__7_ ( .D(n2044), .CK(clk), .RN(rst_n), .Q(
        cal_out[367]) );
  DFFRHQX1 cal_out_reg_11__7_ ( .D(n2284), .CK(clk), .RN(rst_n), .Q(
        cal_out[127]) );
  DFFRHQX1 cal_out_reg_1__8_ ( .D(n1883), .CK(clk), .RN(rst_n), .Q(
        cal_out[528]) );
  DFFRHQX1 cal_out_reg_3__8_ ( .D(n1963), .CK(clk), .RN(rst_n), .Q(
        cal_out[448]) );
  DFFRHQX1 cal_out_reg_5__8_ ( .D(n2043), .CK(clk), .RN(rst_n), .Q(
        cal_out[368]) );
  DFFRHQX1 cal_out_reg_7__8_ ( .D(n2123), .CK(clk), .RN(rst_n), .Q(
        cal_out[288]) );
  DFFRHQX1 cal_out_reg_11__8_ ( .D(n2283), .CK(clk), .RN(rst_n), .Q(
        cal_out[128]) );
  DFFRHQX1 cal_out_reg_13__8_ ( .D(n2363), .CK(clk), .RN(rst_n), .Q(
        cal_out[48]) );
  DFFRHQX1 cal_out_reg_5__9_ ( .D(n2042), .CK(clk), .RN(rst_n), .Q(
        cal_out[369]) );
  DFFRHQX1 cal_out_reg_11__9_ ( .D(n2282), .CK(clk), .RN(rst_n), .Q(
        cal_out[129]) );
  DFFRHQX1 cal_out_reg_5__11_ ( .D(n2040), .CK(clk), .RN(rst_n), .Q(
        cal_out[371]) );
  DFFRHQX1 cal_out_reg_11__11_ ( .D(n2280), .CK(clk), .RN(rst_n), .Q(
        cal_out[131]) );
  DFFRHQX1 cal_out_reg_1__12_ ( .D(n1879), .CK(clk), .RN(rst_n), .Q(
        cal_out[532]) );
  DFFRHQX1 cal_out_reg_3__12_ ( .D(n1959), .CK(clk), .RN(rst_n), .Q(
        cal_out[452]) );
  DFFRHQX1 cal_out_reg_5__12_ ( .D(n2039), .CK(clk), .RN(rst_n), .Q(
        cal_out[372]) );
  DFFRHQX1 cal_out_reg_7__12_ ( .D(n2119), .CK(clk), .RN(rst_n), .Q(
        cal_out[292]) );
  DFFRHQX1 cal_out_reg_11__12_ ( .D(n2279), .CK(clk), .RN(rst_n), .Q(
        cal_out[132]) );
  DFFRHQX1 cal_out_reg_13__12_ ( .D(n2359), .CK(clk), .RN(rst_n), .Q(
        cal_out[52]) );
  DFFRHQX1 cal_out_reg_5__13_ ( .D(n2038), .CK(clk), .RN(rst_n), .Q(
        cal_out[373]) );
  DFFRHQX1 cal_out_reg_7__13_ ( .D(n2118), .CK(clk), .RN(rst_n), .Q(
        cal_out[293]) );
  DFFRHQX1 cal_out_reg_11__13_ ( .D(n2278), .CK(clk), .RN(rst_n), .Q(
        cal_out[133]) );
  DFFRHQX1 cal_out_reg_1__14_ ( .D(n1877), .CK(clk), .RN(rst_n), .Q(
        cal_out[534]) );
  DFFRHQX1 cal_out_reg_3__14_ ( .D(n1957), .CK(clk), .RN(rst_n), .Q(
        cal_out[454]) );
  DFFRHQX1 cal_out_reg_5__14_ ( .D(n2037), .CK(clk), .RN(rst_n), .Q(
        cal_out[374]) );
  DFFRHQX1 cal_out_reg_7__14_ ( .D(n2117), .CK(clk), .RN(rst_n), .Q(
        cal_out[294]) );
  DFFRHQX1 cal_out_reg_11__14_ ( .D(n2277), .CK(clk), .RN(rst_n), .Q(
        cal_out[134]) );
  DFFRHQX1 cal_out_reg_13__14_ ( .D(n2357), .CK(clk), .RN(rst_n), .Q(
        cal_out[54]) );
  DFFRHQX1 cal_out_reg_5__15_ ( .D(n2036), .CK(clk), .RN(rst_n), .Q(
        cal_out[375]) );
  DFFRHQX1 cal_out_reg_7__15_ ( .D(n2116), .CK(clk), .RN(rst_n), .Q(
        cal_out[295]) );
  DFFRHQX1 cal_out_reg_11__15_ ( .D(n2276), .CK(clk), .RN(rst_n), .Q(
        cal_out[135]) );
  DFFRHQX1 cal_out_reg_1__16_ ( .D(n1875), .CK(clk), .RN(rst_n), .Q(
        cal_out[536]) );
  DFFRHQX1 cal_out_reg_3__16_ ( .D(n1955), .CK(clk), .RN(rst_n), .Q(
        cal_out[456]) );
  DFFRHQX1 cal_out_reg_5__16_ ( .D(n2035), .CK(clk), .RN(rst_n), .Q(
        cal_out[376]) );
  DFFRHQX1 cal_out_reg_7__16_ ( .D(n2115), .CK(clk), .RN(rst_n), .Q(
        cal_out[296]) );
  DFFRHQX1 cal_out_reg_11__16_ ( .D(n2275), .CK(clk), .RN(rst_n), .Q(
        cal_out[136]) );
  DFFRHQX1 cal_out_reg_13__16_ ( .D(n2355), .CK(clk), .RN(rst_n), .Q(
        cal_out[56]) );
  DFFRHQX1 cal_out_reg_1__17_ ( .D(n1874), .CK(clk), .RN(rst_n), .Q(
        cal_out[537]) );
  DFFRHQX1 cal_out_reg_3__17_ ( .D(n1954), .CK(clk), .RN(rst_n), .Q(
        cal_out[457]) );
  DFFRHQX1 cal_out_reg_5__17_ ( .D(n2034), .CK(clk), .RN(rst_n), .Q(
        cal_out[377]) );
  DFFRHQX1 cal_out_reg_7__17_ ( .D(n2114), .CK(clk), .RN(rst_n), .Q(
        cal_out[297]) );
  DFFRHQX1 cal_out_reg_11__17_ ( .D(n2274), .CK(clk), .RN(rst_n), .Q(
        cal_out[137]) );
  DFFRHQX1 cal_out_reg_13__17_ ( .D(n2354), .CK(clk), .RN(rst_n), .Q(
        cal_out[57]) );
  DFFRHQX1 cal_out_reg_5__18_ ( .D(n2033), .CK(clk), .RN(rst_n), .Q(
        cal_out[378]) );
  DFFRHQX1 cal_out_reg_11__18_ ( .D(n2273), .CK(clk), .RN(rst_n), .Q(
        cal_out[138]) );
  DFFRHQX1 cal_out_reg_5__19_ ( .D(n2032), .CK(clk), .RN(rst_n), .Q(
        cal_out[379]) );
  DFFRHQX1 cal_out_reg_11__19_ ( .D(n2272), .CK(clk), .RN(rst_n), .Q(
        cal_out[139]) );
  DFFRHQX1 cal_out_reg_1__20_ ( .D(n1871), .CK(clk), .RN(rst_n), .Q(
        cal_out[540]) );
  DFFRHQX1 cal_out_reg_3__20_ ( .D(n1951), .CK(clk), .RN(rst_n), .Q(
        cal_out[460]) );
  DFFRHQX1 cal_out_reg_5__20_ ( .D(n2031), .CK(clk), .RN(rst_n), .Q(
        cal_out[380]) );
  DFFRHQX1 cal_out_reg_7__20_ ( .D(n2111), .CK(clk), .RN(rst_n), .Q(
        cal_out[300]) );
  DFFRHQX1 cal_out_reg_11__20_ ( .D(n2271), .CK(clk), .RN(rst_n), .Q(
        cal_out[140]) );
  DFFRHQX1 cal_out_reg_13__20_ ( .D(n2351), .CK(clk), .RN(rst_n), .Q(
        cal_out[60]) );
  DFFRHQX1 cal_out_reg_1__21_ ( .D(n1870), .CK(clk), .RN(rst_n), .Q(
        cal_out[541]) );
  DFFRHQX1 cal_out_reg_3__21_ ( .D(n1950), .CK(clk), .RN(rst_n), .Q(
        cal_out[461]) );
  DFFRHQX1 cal_out_reg_5__21_ ( .D(n2030), .CK(clk), .RN(rst_n), .Q(
        cal_out[381]) );
  DFFRHQX1 cal_out_reg_7__21_ ( .D(n2110), .CK(clk), .RN(rst_n), .Q(
        cal_out[301]) );
  DFFRHQX1 cal_out_reg_11__21_ ( .D(n2270), .CK(clk), .RN(rst_n), .Q(
        cal_out[141]) );
  DFFRHQX1 cal_out_reg_13__21_ ( .D(n2350), .CK(clk), .RN(rst_n), .Q(
        cal_out[61]) );
  DFFRHQX1 cal_out_reg_1__22_ ( .D(n1869), .CK(clk), .RN(rst_n), .Q(
        cal_out[542]) );
  DFFRHQX1 cal_out_reg_3__22_ ( .D(n1949), .CK(clk), .RN(rst_n), .Q(
        cal_out[462]) );
  DFFRHQX1 cal_out_reg_5__22_ ( .D(n2029), .CK(clk), .RN(rst_n), .Q(
        cal_out[382]) );
  DFFRHQX1 cal_out_reg_7__22_ ( .D(n2109), .CK(clk), .RN(rst_n), .Q(
        cal_out[302]) );
  DFFRHQX1 cal_out_reg_11__22_ ( .D(n2269), .CK(clk), .RN(rst_n), .Q(
        cal_out[142]) );
  DFFRHQX1 cal_out_reg_13__22_ ( .D(n2349), .CK(clk), .RN(rst_n), .Q(
        cal_out[62]) );
  DFFRHQX1 cal_out_reg_1__23_ ( .D(n1868), .CK(clk), .RN(rst_n), .Q(
        cal_out[543]) );
  DFFRHQX1 cal_out_reg_3__23_ ( .D(n1948), .CK(clk), .RN(rst_n), .Q(
        cal_out[463]) );
  DFFRHQX1 cal_out_reg_5__23_ ( .D(n2028), .CK(clk), .RN(rst_n), .Q(
        cal_out[383]) );
  DFFRHQX1 cal_out_reg_7__23_ ( .D(n2108), .CK(clk), .RN(rst_n), .Q(
        cal_out[303]) );
  DFFRHQX1 cal_out_reg_11__23_ ( .D(n2268), .CK(clk), .RN(rst_n), .Q(
        cal_out[143]) );
  DFFRHQX1 cal_out_reg_13__23_ ( .D(n2348), .CK(clk), .RN(rst_n), .Q(
        cal_out[63]) );
  DFFRHQX1 cal_out_reg_1__24_ ( .D(n1867), .CK(clk), .RN(rst_n), .Q(
        cal_out[544]) );
  DFFRHQX1 cal_out_reg_3__24_ ( .D(n1947), .CK(clk), .RN(rst_n), .Q(
        cal_out[464]) );
  DFFRHQX1 cal_out_reg_5__24_ ( .D(n2027), .CK(clk), .RN(rst_n), .Q(
        cal_out[384]) );
  DFFRHQX1 cal_out_reg_7__24_ ( .D(n2107), .CK(clk), .RN(rst_n), .Q(
        cal_out[304]) );
  DFFRHQX1 cal_out_reg_11__24_ ( .D(n2267), .CK(clk), .RN(rst_n), .Q(
        cal_out[144]) );
  DFFRHQX1 cal_out_reg_13__24_ ( .D(n2347), .CK(clk), .RN(rst_n), .Q(
        cal_out[64]) );
  DFFRHQX1 cal_out_reg_1__25_ ( .D(n1866), .CK(clk), .RN(rst_n), .Q(
        cal_out[545]) );
  DFFRHQX1 cal_out_reg_3__25_ ( .D(n1946), .CK(clk), .RN(rst_n), .Q(
        cal_out[465]) );
  DFFRHQX1 cal_out_reg_5__25_ ( .D(n2026), .CK(clk), .RN(rst_n), .Q(
        cal_out[385]) );
  DFFRHQX1 cal_out_reg_7__25_ ( .D(n2106), .CK(clk), .RN(rst_n), .Q(
        cal_out[305]) );
  DFFRHQX1 cal_out_reg_11__25_ ( .D(n2266), .CK(clk), .RN(rst_n), .Q(
        cal_out[145]) );
  DFFRHQX1 cal_out_reg_13__25_ ( .D(n2346), .CK(clk), .RN(rst_n), .Q(
        cal_out[65]) );
  DFFRHQX1 cal_out_reg_5__26_ ( .D(n2025), .CK(clk), .RN(rst_n), .Q(
        cal_out[386]) );
  DFFRHQX1 cal_out_reg_11__26_ ( .D(n2265), .CK(clk), .RN(rst_n), .Q(
        cal_out[146]) );
  DFFRHQX1 cal_out_reg_5__27_ ( .D(n2024), .CK(clk), .RN(rst_n), .Q(
        cal_out[387]) );
  DFFRHQX1 cal_out_reg_11__27_ ( .D(n2264), .CK(clk), .RN(rst_n), .Q(
        cal_out[147]) );
  DFFRHQX1 cal_out_reg_1__28_ ( .D(n1863), .CK(clk), .RN(rst_n), .Q(
        cal_out[548]) );
  DFFRHQX1 cal_out_reg_3__28_ ( .D(n1943), .CK(clk), .RN(rst_n), .Q(
        cal_out[468]) );
  DFFRHQX1 cal_out_reg_5__28_ ( .D(n2023), .CK(clk), .RN(rst_n), .Q(
        cal_out[388]) );
  DFFRHQX1 cal_out_reg_7__28_ ( .D(n2103), .CK(clk), .RN(rst_n), .Q(
        cal_out[308]) );
  DFFRHQX1 cal_out_reg_11__28_ ( .D(n2263), .CK(clk), .RN(rst_n), .Q(
        cal_out[148]) );
  DFFRHQX1 cal_out_reg_13__28_ ( .D(n2343), .CK(clk), .RN(rst_n), .Q(
        cal_out[68]) );
  DFFRHQX1 cal_out_reg_1__29_ ( .D(n1862), .CK(clk), .RN(rst_n), .Q(
        cal_out[549]) );
  DFFRHQX1 cal_out_reg_3__29_ ( .D(n1942), .CK(clk), .RN(rst_n), .Q(
        cal_out[469]) );
  DFFRHQX1 cal_out_reg_5__29_ ( .D(n2022), .CK(clk), .RN(rst_n), .Q(
        cal_out[389]) );
  DFFRHQX1 cal_out_reg_7__29_ ( .D(n2102), .CK(clk), .RN(rst_n), .Q(
        cal_out[309]) );
  DFFRHQX1 cal_out_reg_11__29_ ( .D(n2262), .CK(clk), .RN(rst_n), .Q(
        cal_out[149]) );
  DFFRHQX1 cal_out_reg_13__29_ ( .D(n2342), .CK(clk), .RN(rst_n), .Q(
        cal_out[69]) );
  DFFRHQX1 cal_out_reg_1__30_ ( .D(n1861), .CK(clk), .RN(rst_n), .Q(
        cal_out[550]) );
  DFFRHQX1 cal_out_reg_3__30_ ( .D(n1941), .CK(clk), .RN(rst_n), .Q(
        cal_out[470]) );
  DFFRHQX1 cal_out_reg_5__30_ ( .D(n2021), .CK(clk), .RN(rst_n), .Q(
        cal_out[390]) );
  DFFRHQX1 cal_out_reg_7__30_ ( .D(n2101), .CK(clk), .RN(rst_n), .Q(
        cal_out[310]) );
  DFFRHQX1 cal_out_reg_11__30_ ( .D(n2261), .CK(clk), .RN(rst_n), .Q(
        cal_out[150]) );
  DFFRHQX1 cal_out_reg_13__30_ ( .D(n2341), .CK(clk), .RN(rst_n), .Q(
        cal_out[70]) );
  DFFRHQX1 cal_out_reg_1__31_ ( .D(n1860), .CK(clk), .RN(rst_n), .Q(
        cal_out[551]) );
  DFFRHQX1 cal_out_reg_3__31_ ( .D(n1940), .CK(clk), .RN(rst_n), .Q(
        cal_out[471]) );
  DFFRHQX1 cal_out_reg_5__31_ ( .D(n2020), .CK(clk), .RN(rst_n), .Q(
        cal_out[391]) );
  DFFRHQX1 cal_out_reg_7__31_ ( .D(n2100), .CK(clk), .RN(rst_n), .Q(
        cal_out[311]) );
  DFFRHQX1 cal_out_reg_11__31_ ( .D(n2260), .CK(clk), .RN(rst_n), .Q(
        cal_out[151]) );
  DFFRHQX1 cal_out_reg_13__31_ ( .D(n2340), .CK(clk), .RN(rst_n), .Q(
        cal_out[71]) );
  DFFRHQX1 cal_out_reg_1__32_ ( .D(n1859), .CK(clk), .RN(rst_n), .Q(
        cal_out[552]) );
  DFFRHQX1 cal_out_reg_3__32_ ( .D(n1939), .CK(clk), .RN(rst_n), .Q(
        cal_out[472]) );
  DFFRHQX1 cal_out_reg_7__32_ ( .D(n2099), .CK(clk), .RN(rst_n), .Q(
        cal_out[312]) );
  DFFRHQX1 cal_out_reg_13__32_ ( .D(n2339), .CK(clk), .RN(rst_n), .Q(
        cal_out[72]) );
  DFFRHQX1 cal_out_reg_1__33_ ( .D(n1858), .CK(clk), .RN(rst_n), .Q(
        cal_out[553]) );
  DFFRHQX1 cal_out_reg_3__33_ ( .D(n1938), .CK(clk), .RN(rst_n), .Q(
        cal_out[473]) );
  DFFRHQX1 cal_out_reg_5__33_ ( .D(n2018), .CK(clk), .RN(rst_n), .Q(
        cal_out[393]) );
  DFFRHQX1 cal_out_reg_7__33_ ( .D(n2098), .CK(clk), .RN(rst_n), .Q(
        cal_out[313]) );
  DFFRHQX1 cal_out_reg_11__33_ ( .D(n2258), .CK(clk), .RN(rst_n), .Q(
        cal_out[153]) );
  DFFRHQX1 cal_out_reg_13__33_ ( .D(n2338), .CK(clk), .RN(rst_n), .Q(
        cal_out[73]) );
  DFFRHQX1 cal_out_reg_1__34_ ( .D(n1857), .CK(clk), .RN(rst_n), .Q(
        cal_out[554]) );
  DFFRHQX1 cal_out_reg_3__34_ ( .D(n1937), .CK(clk), .RN(rst_n), .Q(
        cal_out[474]) );
  DFFRHQX1 cal_out_reg_5__34_ ( .D(n2017), .CK(clk), .RN(rst_n), .Q(
        cal_out[394]) );
  DFFRHQX1 cal_out_reg_7__34_ ( .D(n2097), .CK(clk), .RN(rst_n), .Q(
        cal_out[314]) );
  DFFRHQX1 cal_out_reg_11__34_ ( .D(n2257), .CK(clk), .RN(rst_n), .Q(
        cal_out[154]) );
  DFFRHQX1 cal_out_reg_13__34_ ( .D(n2337), .CK(clk), .RN(rst_n), .Q(
        cal_out[74]) );
  DFFRHQX1 cal_out_reg_1__35_ ( .D(n1856), .CK(clk), .RN(rst_n), .Q(
        cal_out[555]) );
  DFFRHQX1 cal_out_reg_3__35_ ( .D(n1936), .CK(clk), .RN(rst_n), .Q(
        cal_out[475]) );
  DFFRHQX1 cal_out_reg_5__35_ ( .D(n2016), .CK(clk), .RN(rst_n), .Q(
        cal_out[395]) );
  DFFRHQX1 cal_out_reg_7__35_ ( .D(n2096), .CK(clk), .RN(rst_n), .Q(
        cal_out[315]) );
  DFFRHQX1 cal_out_reg_11__35_ ( .D(n2256), .CK(clk), .RN(rst_n), .Q(
        cal_out[155]) );
  DFFRHQX1 cal_out_reg_13__35_ ( .D(n2336), .CK(clk), .RN(rst_n), .Q(
        cal_out[75]) );
  DFFRHQX1 cal_out_reg_1__36_ ( .D(n1855), .CK(clk), .RN(rst_n), .Q(
        cal_out[556]) );
  DFFRHQX1 cal_out_reg_3__36_ ( .D(n1935), .CK(clk), .RN(rst_n), .Q(
        cal_out[476]) );
  DFFRHQX1 cal_out_reg_5__36_ ( .D(n2015), .CK(clk), .RN(rst_n), .Q(
        cal_out[396]) );
  DFFRHQX1 cal_out_reg_7__36_ ( .D(n2095), .CK(clk), .RN(rst_n), .Q(
        cal_out[316]) );
  DFFRHQX1 cal_out_reg_11__36_ ( .D(n2255), .CK(clk), .RN(rst_n), .Q(
        cal_out[156]) );
  DFFRHQX1 cal_out_reg_13__36_ ( .D(n2335), .CK(clk), .RN(rst_n), .Q(
        cal_out[76]) );
  DFFRHQX1 cal_out_reg_1__37_ ( .D(n1854), .CK(clk), .RN(rst_n), .Q(
        cal_out[557]) );
  DFFRHQX1 cal_out_reg_3__37_ ( .D(n1934), .CK(clk), .RN(rst_n), .Q(
        cal_out[477]) );
  DFFRHQX1 cal_out_reg_5__37_ ( .D(n2014), .CK(clk), .RN(rst_n), .Q(
        cal_out[397]) );
  DFFRHQX1 cal_out_reg_7__37_ ( .D(n2094), .CK(clk), .RN(rst_n), .Q(
        cal_out[317]) );
  DFFRHQX1 cal_out_reg_11__37_ ( .D(n2254), .CK(clk), .RN(rst_n), .Q(
        cal_out[157]) );
  DFFRHQX1 cal_out_reg_13__37_ ( .D(n2334), .CK(clk), .RN(rst_n), .Q(
        cal_out[77]) );
  DFFRHQX1 cal_out_reg_1__38_ ( .D(n1853), .CK(clk), .RN(rst_n), .Q(
        cal_out[558]) );
  DFFRHQX1 cal_out_reg_3__38_ ( .D(n1933), .CK(clk), .RN(rst_n), .Q(
        cal_out[478]) );
  DFFRHQX1 cal_out_reg_5__38_ ( .D(n2013), .CK(clk), .RN(rst_n), .Q(
        cal_out[398]) );
  DFFRHQX1 cal_out_reg_7__38_ ( .D(n2093), .CK(clk), .RN(rst_n), .Q(
        cal_out[318]) );
  DFFRHQX1 cal_out_reg_11__38_ ( .D(n2253), .CK(clk), .RN(rst_n), .Q(
        cal_out[158]) );
  DFFRHQX1 cal_out_reg_13__38_ ( .D(n2333), .CK(clk), .RN(rst_n), .Q(
        cal_out[78]) );
  DFFRHQX1 cal_out_reg_1__39_ ( .D(n1852), .CK(clk), .RN(rst_n), .Q(
        cal_out[559]) );
  DFFRHQX1 cal_out_reg_3__39_ ( .D(n1932), .CK(clk), .RN(rst_n), .Q(
        cal_out[479]) );
  DFFRHQX1 cal_out_reg_5__39_ ( .D(n2012), .CK(clk), .RN(rst_n), .Q(
        cal_out[399]) );
  DFFRHQX1 cal_out_reg_7__39_ ( .D(n2092), .CK(clk), .RN(rst_n), .Q(
        cal_out[319]) );
  DFFRHQX1 cal_out_reg_11__39_ ( .D(n2252), .CK(clk), .RN(rst_n), .Q(
        cal_out[159]) );
  DFFRHQX1 cal_out_reg_13__39_ ( .D(n2332), .CK(clk), .RN(rst_n), .Q(
        cal_out[79]) );
  DFFRHQX1 length_reg_reg_1__5_ ( .D(n1728), .CK(clk), .RN(rst_n), .Q(
        length_reg[83]) );
  DFFRHQX1 length_reg_reg_3__5_ ( .D(n1740), .CK(clk), .RN(rst_n), .Q(
        length_reg[71]) );
  DFFRHQX1 length_reg_reg_5__5_ ( .D(n1752), .CK(clk), .RN(rst_n), .Q(
        length_reg[59]) );
  DFFRHQX1 length_reg_reg_7__5_ ( .D(n1764), .CK(clk), .RN(rst_n), .Q(
        length_reg[47]) );
  DFFRHQX1 length_reg_reg_11__5_ ( .D(n1788), .CK(clk), .RN(rst_n), .Q(
        length_reg[23]) );
  DFFRHQX1 length_reg_reg_13__5_ ( .D(n1800), .CK(clk), .RN(rst_n), .Q(
        length_reg[11]) );
  DFFRHQX1 length_reg_reg_1__3_ ( .D(n1730), .CK(clk), .RN(rst_n), .Q(
        length_reg[81]) );
  DFFRHQX1 length_reg_reg_3__3_ ( .D(n1742), .CK(clk), .RN(rst_n), .Q(
        length_reg[69]) );
  DFFRHQX1 length_reg_reg_5__3_ ( .D(n1754), .CK(clk), .RN(rst_n), .Q(
        length_reg[57]) );
  DFFRHQX1 length_reg_reg_7__3_ ( .D(n1766), .CK(clk), .RN(rst_n), .Q(
        length_reg[45]) );
  DFFRHQX1 length_reg_reg_11__3_ ( .D(n1790), .CK(clk), .RN(rst_n), .Q(
        length_reg[21]) );
  DFFRHQX1 length_reg_reg_13__3_ ( .D(n1802), .CK(clk), .RN(rst_n), .Q(
        length_reg[9]) );
  DFFRHQX1 length_reg_reg_1__1_ ( .D(n1732), .CK(clk), .RN(rst_n), .Q(
        length_reg[79]) );
  DFFRHQX1 length_reg_reg_3__1_ ( .D(n1744), .CK(clk), .RN(rst_n), .Q(
        length_reg[67]) );
  DFFRHQX1 length_reg_reg_5__1_ ( .D(n1756), .CK(clk), .RN(rst_n), .Q(
        length_reg[55]) );
  DFFRHQX1 length_reg_reg_7__1_ ( .D(n1768), .CK(clk), .RN(rst_n), .Q(
        length_reg[43]) );
  DFFRHQX1 length_reg_reg_11__1_ ( .D(n1792), .CK(clk), .RN(rst_n), .Q(
        length_reg[19]) );
  DFFRHQX1 length_reg_reg_13__1_ ( .D(n1804), .CK(clk), .RN(rst_n), .Q(
        length_reg[7]) );
  DFFRHQX1 length_reg_reg_1__4_ ( .D(n1729), .CK(clk), .RN(rst_n), .Q(
        length_reg[82]) );
  DFFRHQX1 length_reg_reg_3__4_ ( .D(n1741), .CK(clk), .RN(rst_n), .Q(
        length_reg[70]) );
  DFFRHQX1 length_reg_reg_5__4_ ( .D(n1753), .CK(clk), .RN(rst_n), .Q(
        length_reg[58]) );
  DFFRHQX1 length_reg_reg_7__4_ ( .D(n1765), .CK(clk), .RN(rst_n), .Q(
        length_reg[46]) );
  DFFRHQX1 length_reg_reg_11__4_ ( .D(n1789), .CK(clk), .RN(rst_n), .Q(
        length_reg[22]) );
  DFFRHQX1 length_reg_reg_13__4_ ( .D(n1801), .CK(clk), .RN(rst_n), .Q(
        length_reg[10]) );
  DFFRHQX1 length_reg_reg_1__2_ ( .D(n1731), .CK(clk), .RN(rst_n), .Q(
        length_reg[80]) );
  DFFRHQX1 length_reg_reg_3__2_ ( .D(n1743), .CK(clk), .RN(rst_n), .Q(
        length_reg[68]) );
  DFFRHQX1 length_reg_reg_5__2_ ( .D(n1755), .CK(clk), .RN(rst_n), .Q(
        length_reg[56]) );
  DFFRHQX1 length_reg_reg_7__2_ ( .D(n1767), .CK(clk), .RN(rst_n), .Q(
        length_reg[44]) );
  DFFRHQX1 length_reg_reg_11__2_ ( .D(n1791), .CK(clk), .RN(rst_n), .Q(
        length_reg[20]) );
  DFFRHQX1 length_reg_reg_13__2_ ( .D(n1803), .CK(clk), .RN(rst_n), .Q(
        length_reg[8]) );
  DFFRHQX1 length_reg_reg_1__0_ ( .D(n1733), .CK(clk), .RN(rst_n), .Q(
        length_reg[78]) );
  DFFRHQX1 length_reg_reg_5__0_ ( .D(n1757), .CK(clk), .RN(rst_n), .Q(
        length_reg[54]) );
  DFFRHQX1 length_reg_reg_7__0_ ( .D(n1769), .CK(clk), .RN(rst_n), .Q(
        length_reg[42]) );
  DFFRHQX1 length_reg_reg_11__0_ ( .D(n1793), .CK(clk), .RN(rst_n), .Q(
        length_reg[18]) );
  DFFRHQX1 cal_out_reg_9__0_ ( .D(n2211), .CK(clk), .RN(rst_n), .Q(
        cal_out[200]) );
  DFFRHQX1 cal_out_reg_9__4_ ( .D(n2207), .CK(clk), .RN(rst_n), .Q(
        cal_out[204]) );
  DFFRHQX1 cal_out_reg_9__5_ ( .D(n2206), .CK(clk), .RN(rst_n), .Q(
        cal_out[205]) );
  DFFRHQX1 cal_out_reg_9__6_ ( .D(n2205), .CK(clk), .RN(rst_n), .Q(
        cal_out[206]) );
  DFFRHQX1 cal_out_reg_9__7_ ( .D(n2204), .CK(clk), .RN(rst_n), .Q(
        cal_out[207]) );
  DFFRHQX1 cal_out_reg_9__8_ ( .D(n2203), .CK(clk), .RN(rst_n), .Q(
        cal_out[208]) );
  DFFRHQX1 cal_out_reg_9__12_ ( .D(n2199), .CK(clk), .RN(rst_n), .Q(
        cal_out[212]) );
  DFFRHQX1 cal_out_reg_9__13_ ( .D(n2198), .CK(clk), .RN(rst_n), .Q(
        cal_out[213]) );
  DFFRHQX1 cal_out_reg_9__14_ ( .D(n2197), .CK(clk), .RN(rst_n), .Q(
        cal_out[214]) );
  DFFRHQX1 cal_out_reg_9__15_ ( .D(n2196), .CK(clk), .RN(rst_n), .Q(
        cal_out[215]) );
  DFFRHQX1 cal_out_reg_9__16_ ( .D(n2195), .CK(clk), .RN(rst_n), .Q(
        cal_out[216]) );
  DFFRHQX1 cal_out_reg_9__17_ ( .D(n2194), .CK(clk), .RN(rst_n), .Q(
        cal_out[217]) );
  DFFRHQX1 cal_out_reg_9__20_ ( .D(n2191), .CK(clk), .RN(rst_n), .Q(
        cal_out[220]) );
  DFFRHQX1 cal_out_reg_9__21_ ( .D(n2190), .CK(clk), .RN(rst_n), .Q(
        cal_out[221]) );
  DFFRHQX1 cal_out_reg_9__22_ ( .D(n2189), .CK(clk), .RN(rst_n), .Q(
        cal_out[222]) );
  DFFRHQX1 cal_out_reg_9__23_ ( .D(n2188), .CK(clk), .RN(rst_n), .Q(
        cal_out[223]) );
  DFFRHQX1 cal_out_reg_9__24_ ( .D(n2187), .CK(clk), .RN(rst_n), .Q(
        cal_out[224]) );
  DFFRHQX1 cal_out_reg_9__25_ ( .D(n2186), .CK(clk), .RN(rst_n), .Q(
        cal_out[225]) );
  DFFRHQX1 cal_out_reg_9__28_ ( .D(n2183), .CK(clk), .RN(rst_n), .Q(
        cal_out[228]) );
  DFFRHQX1 cal_out_reg_9__29_ ( .D(n2182), .CK(clk), .RN(rst_n), .Q(
        cal_out[229]) );
  DFFRHQX1 cal_out_reg_9__30_ ( .D(n2181), .CK(clk), .RN(rst_n), .Q(
        cal_out[230]) );
  DFFRHQX1 cal_out_reg_9__31_ ( .D(n2180), .CK(clk), .RN(rst_n), .Q(
        cal_out[231]) );
  DFFRHQX1 cal_out_reg_9__32_ ( .D(n2179), .CK(clk), .RN(rst_n), .Q(
        cal_out[232]) );
  DFFRHQX1 cal_out_reg_9__33_ ( .D(n2178), .CK(clk), .RN(rst_n), .Q(
        cal_out[233]) );
  DFFRHQX1 cal_out_reg_9__34_ ( .D(n2177), .CK(clk), .RN(rst_n), .Q(
        cal_out[234]) );
  DFFRHQX1 cal_out_reg_9__35_ ( .D(n2176), .CK(clk), .RN(rst_n), .Q(
        cal_out[235]) );
  DFFRHQX1 cal_out_reg_9__36_ ( .D(n2175), .CK(clk), .RN(rst_n), .Q(
        cal_out[236]) );
  DFFRHQX1 cal_out_reg_9__37_ ( .D(n2174), .CK(clk), .RN(rst_n), .Q(
        cal_out[237]) );
  DFFRHQX1 cal_out_reg_9__38_ ( .D(n2173), .CK(clk), .RN(rst_n), .Q(
        cal_out[238]) );
  DFFRHQX1 cal_out_reg_9__39_ ( .D(n2172), .CK(clk), .RN(rst_n), .Q(
        cal_out[239]) );
  DFFRHQX1 length_reg_reg_9__5_ ( .D(n1776), .CK(clk), .RN(rst_n), .Q(
        length_reg[35]) );
  DFFRHQX1 length_reg_reg_9__3_ ( .D(n1778), .CK(clk), .RN(rst_n), .Q(
        length_reg[33]) );
  DFFRHQX1 length_reg_reg_9__1_ ( .D(n1780), .CK(clk), .RN(rst_n), .Q(
        length_reg[31]) );
  DFFRHQX1 length_reg_reg_9__4_ ( .D(n1777), .CK(clk), .RN(rst_n), .Q(
        length_reg[34]) );
  DFFRHQX1 length_reg_reg_9__2_ ( .D(n1779), .CK(clk), .RN(rst_n), .Q(
        length_reg[32]) );
  DFFRHQX1 length_reg_reg_9__0_ ( .D(n1781), .CK(clk), .RN(rst_n), .Q(
        length_reg[30]) );
  DFFRHQX1 cal_out_reg_8__0_ ( .D(n2171), .CK(clk), .RN(rst_n), .Q(
        cal_out[240]) );
  DFFRHQX1 cal_out_reg_8__1_ ( .D(n2170), .CK(clk), .RN(rst_n), .Q(
        cal_out[241]) );
  DFFRHQX1 cal_out_reg_8__4_ ( .D(n2167), .CK(clk), .RN(rst_n), .Q(
        cal_out[244]) );
  DFFRHQX1 cal_out_reg_8__5_ ( .D(n2166), .CK(clk), .RN(rst_n), .Q(
        cal_out[245]) );
  DFFRHQX1 cal_out_reg_8__6_ ( .D(n2165), .CK(clk), .RN(rst_n), .Q(
        cal_out[246]) );
  DFFRHQX1 cal_out_reg_8__7_ ( .D(n2164), .CK(clk), .RN(rst_n), .Q(
        cal_out[247]) );
  DFFRHQX1 cal_out_reg_8__8_ ( .D(n2163), .CK(clk), .RN(rst_n), .Q(
        cal_out[248]) );
  DFFRHQX1 cal_out_reg_8__9_ ( .D(n2162), .CK(clk), .RN(rst_n), .Q(
        cal_out[249]) );
  DFFRHQX1 cal_out_reg_8__12_ ( .D(n2159), .CK(clk), .RN(rst_n), .Q(
        cal_out[252]) );
  DFFRHQX1 cal_out_reg_8__13_ ( .D(n2158), .CK(clk), .RN(rst_n), .Q(
        cal_out[253]) );
  DFFRHQX1 cal_out_reg_8__14_ ( .D(n2157), .CK(clk), .RN(rst_n), .Q(
        cal_out[254]) );
  DFFRHQX1 cal_out_reg_8__15_ ( .D(n2156), .CK(clk), .RN(rst_n), .Q(
        cal_out[255]) );
  DFFRHQX1 cal_out_reg_8__16_ ( .D(n2155), .CK(clk), .RN(rst_n), .Q(
        cal_out[256]) );
  DFFRHQX1 cal_out_reg_8__17_ ( .D(n2154), .CK(clk), .RN(rst_n), .Q(
        cal_out[257]) );
  DFFRHQX1 cal_out_reg_8__20_ ( .D(n2151), .CK(clk), .RN(rst_n), .Q(
        cal_out[260]) );
  DFFRHQX1 cal_out_reg_8__21_ ( .D(n2150), .CK(clk), .RN(rst_n), .Q(
        cal_out[261]) );
  DFFRHQX1 cal_out_reg_8__22_ ( .D(n2149), .CK(clk), .RN(rst_n), .Q(
        cal_out[262]) );
  DFFRHQX1 cal_out_reg_8__23_ ( .D(n2148), .CK(clk), .RN(rst_n), .Q(
        cal_out[263]) );
  DFFRHQX1 cal_out_reg_8__24_ ( .D(n2147), .CK(clk), .RN(rst_n), .Q(
        cal_out[264]) );
  DFFRHQX1 cal_out_reg_8__25_ ( .D(n2146), .CK(clk), .RN(rst_n), .Q(
        cal_out[265]) );
  DFFRHQX1 cal_out_reg_8__28_ ( .D(n2143), .CK(clk), .RN(rst_n), .Q(
        cal_out[268]) );
  DFFRHQX1 cal_out_reg_8__29_ ( .D(n2142), .CK(clk), .RN(rst_n), .Q(
        cal_out[269]) );
  DFFRHQX1 cal_out_reg_8__30_ ( .D(n2141), .CK(clk), .RN(rst_n), .Q(
        cal_out[270]) );
  DFFRHQX1 cal_out_reg_8__31_ ( .D(n2140), .CK(clk), .RN(rst_n), .Q(
        cal_out[271]) );
  DFFRHQX1 cal_out_reg_8__32_ ( .D(n2139), .CK(clk), .RN(rst_n), .Q(
        cal_out[272]) );
  DFFRHQX1 cal_out_reg_8__33_ ( .D(n2138), .CK(clk), .RN(rst_n), .Q(
        cal_out[273]) );
  DFFRHQX1 cal_out_reg_8__34_ ( .D(n2137), .CK(clk), .RN(rst_n), .Q(
        cal_out[274]) );
  DFFRHQX1 cal_out_reg_8__35_ ( .D(n2136), .CK(clk), .RN(rst_n), .Q(
        cal_out[275]) );
  DFFRHQX1 cal_out_reg_8__36_ ( .D(n2135), .CK(clk), .RN(rst_n), .Q(
        cal_out[276]) );
  DFFRHQX1 cal_out_reg_8__37_ ( .D(n2134), .CK(clk), .RN(rst_n), .Q(
        cal_out[277]) );
  DFFRHQX1 cal_out_reg_8__38_ ( .D(n2133), .CK(clk), .RN(rst_n), .Q(
        cal_out[278]) );
  DFFRHQX1 cal_out_reg_8__39_ ( .D(n2132), .CK(clk), .RN(rst_n), .Q(
        cal_out[279]) );
  DFFRHQX1 length_reg_reg_8__5_ ( .D(n1770), .CK(clk), .RN(rst_n), .Q(
        length_reg[41]) );
  DFFRHQX1 length_reg_reg_8__3_ ( .D(n1772), .CK(clk), .RN(rst_n), .Q(
        length_reg[39]) );
  DFFRHQX1 length_reg_reg_8__1_ ( .D(n1774), .CK(clk), .RN(rst_n), .Q(
        length_reg[37]) );
  DFFRHQX1 length_reg_reg_8__4_ ( .D(n1771), .CK(clk), .RN(rst_n), .Q(
        length_reg[40]) );
  DFFRHQX1 length_reg_reg_8__2_ ( .D(n1773), .CK(clk), .RN(rst_n), .Q(
        length_reg[38]) );
  DFFRHQX1 length_reg_reg_8__0_ ( .D(n1775), .CK(clk), .RN(rst_n), .Q(
        length_reg[36]) );
  DFFRHQX1 cal_out_reg_0__0_ ( .D(n1851), .CK(clk), .RN(rst_n), .Q(
        cal_out[560]) );
  DFFRHQX1 cal_out_reg_2__0_ ( .D(n1931), .CK(clk), .RN(rst_n), .Q(
        cal_out[480]) );
  DFFRHQX1 cal_out_reg_4__0_ ( .D(n2011), .CK(clk), .RN(rst_n), .Q(
        cal_out[400]) );
  DFFRHQX1 cal_out_reg_6__0_ ( .D(n2091), .CK(clk), .RN(rst_n), .Q(
        cal_out[320]) );
  DFFRHQX1 cal_out_reg_12__0_ ( .D(n2331), .CK(clk), .RN(rst_n), .Q(
        cal_out[80]) );
  DFFRHQX1 cal_out_reg_14__0_ ( .D(n2411), .CK(clk), .RN(rst_n), .Q(cal_out[0]) );
  DFFRHQX1 cal_out_reg_2__1_ ( .D(n1930), .CK(clk), .RN(rst_n), .Q(
        cal_out[481]) );
  DFFRHQX1 cal_out_reg_4__1_ ( .D(n2010), .CK(clk), .RN(rst_n), .Q(
        cal_out[401]) );
  DFFRHQX1 cal_out_reg_6__1_ ( .D(n2090), .CK(clk), .RN(rst_n), .Q(
        cal_out[321]) );
  DFFRHQX1 cal_out_reg_4__2_ ( .D(n2009), .CK(clk), .RN(rst_n), .Q(
        cal_out[402]) );
  DFFRHQX1 cal_out_reg_6__2_ ( .D(n2089), .CK(clk), .RN(rst_n), .Q(
        cal_out[322]) );
  DFFRHQX1 cal_out_reg_4__3_ ( .D(n2008), .CK(clk), .RN(rst_n), .Q(
        cal_out[403]) );
  DFFRHQX1 cal_out_reg_6__3_ ( .D(n2088), .CK(clk), .RN(rst_n), .Q(
        cal_out[323]) );
  DFFRHQX1 cal_out_reg_0__4_ ( .D(n1847), .CK(clk), .RN(rst_n), .Q(
        cal_out[564]) );
  DFFRHQX1 cal_out_reg_2__4_ ( .D(n1927), .CK(clk), .RN(rst_n), .Q(
        cal_out[484]) );
  DFFRHQX1 cal_out_reg_4__4_ ( .D(n2007), .CK(clk), .RN(rst_n), .Q(
        cal_out[404]) );
  DFFRHQX1 cal_out_reg_6__4_ ( .D(n2087), .CK(clk), .RN(rst_n), .Q(
        cal_out[324]) );
  DFFRHQX1 cal_out_reg_12__4_ ( .D(n2327), .CK(clk), .RN(rst_n), .Q(
        cal_out[84]) );
  DFFRHQX1 cal_out_reg_14__4_ ( .D(n2407), .CK(clk), .RN(rst_n), .Q(cal_out[4]) );
  DFFRHQX1 cal_out_reg_0__5_ ( .D(n1846), .CK(clk), .RN(rst_n), .Q(
        cal_out[565]) );
  DFFRHQX1 cal_out_reg_2__5_ ( .D(n1926), .CK(clk), .RN(rst_n), .Q(
        cal_out[485]) );
  DFFRHQX1 cal_out_reg_4__5_ ( .D(n2006), .CK(clk), .RN(rst_n), .Q(
        cal_out[405]) );
  DFFRHQX1 cal_out_reg_6__5_ ( .D(n2086), .CK(clk), .RN(rst_n), .Q(
        cal_out[325]) );
  DFFRHQX1 cal_out_reg_12__5_ ( .D(n2326), .CK(clk), .RN(rst_n), .Q(
        cal_out[85]) );
  DFFRHQX1 cal_out_reg_14__5_ ( .D(n2406), .CK(clk), .RN(rst_n), .Q(cal_out[5]) );
  DFFRHQX1 cal_out_reg_0__6_ ( .D(n1845), .CK(clk), .RN(rst_n), .Q(
        cal_out[566]) );
  DFFRHQX1 cal_out_reg_2__6_ ( .D(n1925), .CK(clk), .RN(rst_n), .Q(
        cal_out[486]) );
  DFFRHQX1 cal_out_reg_4__6_ ( .D(n2005), .CK(clk), .RN(rst_n), .Q(
        cal_out[406]) );
  DFFRHQX1 cal_out_reg_6__6_ ( .D(n2085), .CK(clk), .RN(rst_n), .Q(
        cal_out[326]) );
  DFFRHQX1 cal_out_reg_12__6_ ( .D(n2325), .CK(clk), .RN(rst_n), .Q(
        cal_out[86]) );
  DFFRHQX1 cal_out_reg_14__6_ ( .D(n2405), .CK(clk), .RN(rst_n), .Q(cal_out[6]) );
  DFFRHQX1 cal_out_reg_0__7_ ( .D(n1844), .CK(clk), .RN(rst_n), .Q(
        cal_out[567]) );
  DFFRHQX1 cal_out_reg_2__7_ ( .D(n1924), .CK(clk), .RN(rst_n), .Q(
        cal_out[487]) );
  DFFRHQX1 cal_out_reg_4__7_ ( .D(n2004), .CK(clk), .RN(rst_n), .Q(
        cal_out[407]) );
  DFFRHQX1 cal_out_reg_6__7_ ( .D(n2084), .CK(clk), .RN(rst_n), .Q(
        cal_out[327]) );
  DFFRHQX1 cal_out_reg_12__7_ ( .D(n2324), .CK(clk), .RN(rst_n), .Q(
        cal_out[87]) );
  DFFRHQX1 cal_out_reg_14__7_ ( .D(n2404), .CK(clk), .RN(rst_n), .Q(cal_out[7]) );
  DFFRHQX1 cal_out_reg_0__8_ ( .D(n1843), .CK(clk), .RN(rst_n), .Q(
        cal_out[568]) );
  DFFRHQX1 cal_out_reg_2__8_ ( .D(n1923), .CK(clk), .RN(rst_n), .Q(
        cal_out[488]) );
  DFFRHQX1 cal_out_reg_4__8_ ( .D(n2003), .CK(clk), .RN(rst_n), .Q(
        cal_out[408]) );
  DFFRHQX1 cal_out_reg_6__8_ ( .D(n2083), .CK(clk), .RN(rst_n), .Q(
        cal_out[328]) );
  DFFRHQX1 cal_out_reg_12__8_ ( .D(n2323), .CK(clk), .RN(rst_n), .Q(
        cal_out[88]) );
  DFFRHQX1 cal_out_reg_14__8_ ( .D(n2403), .CK(clk), .RN(rst_n), .Q(cal_out[8]) );
  DFFRHQX1 cal_out_reg_0__9_ ( .D(n1842), .CK(clk), .RN(rst_n), .Q(
        cal_out[569]) );
  DFFRHQX1 cal_out_reg_2__9_ ( .D(n1922), .CK(clk), .RN(rst_n), .Q(
        cal_out[489]) );
  DFFRHQX1 cal_out_reg_4__9_ ( .D(n2002), .CK(clk), .RN(rst_n), .Q(
        cal_out[409]) );
  DFFRHQX1 cal_out_reg_6__9_ ( .D(n2082), .CK(clk), .RN(rst_n), .Q(
        cal_out[329]) );
  DFFRHQX1 cal_out_reg_4__10_ ( .D(n2001), .CK(clk), .RN(rst_n), .Q(
        cal_out[410]) );
  DFFRHQX1 cal_out_reg_6__10_ ( .D(n2081), .CK(clk), .RN(rst_n), .Q(
        cal_out[330]) );
  DFFRHQX1 cal_out_reg_4__11_ ( .D(n2000), .CK(clk), .RN(rst_n), .Q(
        cal_out[411]) );
  DFFRHQX1 cal_out_reg_6__11_ ( .D(n2080), .CK(clk), .RN(rst_n), .Q(
        cal_out[331]) );
  DFFRHQX1 cal_out_reg_0__12_ ( .D(n1839), .CK(clk), .RN(rst_n), .Q(
        cal_out[572]) );
  DFFRHQX1 cal_out_reg_2__12_ ( .D(n1919), .CK(clk), .RN(rst_n), .Q(
        cal_out[492]) );
  DFFRHQX1 cal_out_reg_4__12_ ( .D(n1999), .CK(clk), .RN(rst_n), .Q(
        cal_out[412]) );
  DFFRHQX1 cal_out_reg_6__12_ ( .D(n2079), .CK(clk), .RN(rst_n), .Q(
        cal_out[332]) );
  DFFRHQX1 cal_out_reg_12__12_ ( .D(n2319), .CK(clk), .RN(rst_n), .Q(
        cal_out[92]) );
  DFFRHQX1 cal_out_reg_14__12_ ( .D(n2399), .CK(clk), .RN(rst_n), .Q(
        cal_out[12]) );
  DFFRHQX1 cal_out_reg_0__13_ ( .D(n1838), .CK(clk), .RN(rst_n), .Q(
        cal_out[573]) );
  DFFRHQX1 cal_out_reg_2__13_ ( .D(n1918), .CK(clk), .RN(rst_n), .Q(
        cal_out[493]) );
  DFFRHQX1 cal_out_reg_4__13_ ( .D(n1998), .CK(clk), .RN(rst_n), .Q(
        cal_out[413]) );
  DFFRHQX1 cal_out_reg_6__13_ ( .D(n2078), .CK(clk), .RN(rst_n), .Q(
        cal_out[333]) );
  DFFRHQX1 cal_out_reg_12__13_ ( .D(n2318), .CK(clk), .RN(rst_n), .Q(
        cal_out[93]) );
  DFFRHQX1 cal_out_reg_14__13_ ( .D(n2398), .CK(clk), .RN(rst_n), .Q(
        cal_out[13]) );
  DFFRHQX1 cal_out_reg_0__14_ ( .D(n1837), .CK(clk), .RN(rst_n), .Q(
        cal_out[574]) );
  DFFRHQX1 cal_out_reg_2__14_ ( .D(n1917), .CK(clk), .RN(rst_n), .Q(
        cal_out[494]) );
  DFFRHQX1 cal_out_reg_4__14_ ( .D(n1997), .CK(clk), .RN(rst_n), .Q(
        cal_out[414]) );
  DFFRHQX1 cal_out_reg_6__14_ ( .D(n2077), .CK(clk), .RN(rst_n), .Q(
        cal_out[334]) );
  DFFRHQX1 cal_out_reg_12__14_ ( .D(n2317), .CK(clk), .RN(rst_n), .Q(
        cal_out[94]) );
  DFFRHQX1 cal_out_reg_14__14_ ( .D(n2397), .CK(clk), .RN(rst_n), .Q(
        cal_out[14]) );
  DFFRHQX1 cal_out_reg_0__15_ ( .D(n1836), .CK(clk), .RN(rst_n), .Q(
        cal_out[575]) );
  DFFRHQX1 cal_out_reg_2__15_ ( .D(n1916), .CK(clk), .RN(rst_n), .Q(
        cal_out[495]) );
  DFFRHQX1 cal_out_reg_4__15_ ( .D(n1996), .CK(clk), .RN(rst_n), .Q(
        cal_out[415]) );
  DFFRHQX1 cal_out_reg_6__15_ ( .D(n2076), .CK(clk), .RN(rst_n), .Q(
        cal_out[335]) );
  DFFRHQX1 cal_out_reg_12__15_ ( .D(n2316), .CK(clk), .RN(rst_n), .Q(
        cal_out[95]) );
  DFFRHQX1 cal_out_reg_14__15_ ( .D(n2396), .CK(clk), .RN(rst_n), .Q(
        cal_out[15]) );
  DFFRHQX1 cal_out_reg_0__16_ ( .D(n1835), .CK(clk), .RN(rst_n), .Q(
        cal_out[576]) );
  DFFRHQX1 cal_out_reg_2__16_ ( .D(n1915), .CK(clk), .RN(rst_n), .Q(
        cal_out[496]) );
  DFFRHQX1 cal_out_reg_4__16_ ( .D(n1995), .CK(clk), .RN(rst_n), .Q(
        cal_out[416]) );
  DFFRHQX1 cal_out_reg_6__16_ ( .D(n2075), .CK(clk), .RN(rst_n), .Q(
        cal_out[336]) );
  DFFRHQX1 cal_out_reg_12__16_ ( .D(n2315), .CK(clk), .RN(rst_n), .Q(
        cal_out[96]) );
  DFFRHQX1 cal_out_reg_14__16_ ( .D(n2395), .CK(clk), .RN(rst_n), .Q(
        cal_out[16]) );
  DFFRHQX1 cal_out_reg_0__17_ ( .D(n1834), .CK(clk), .RN(rst_n), .Q(
        cal_out[577]) );
  DFFRHQX1 cal_out_reg_2__17_ ( .D(n1914), .CK(clk), .RN(rst_n), .Q(
        cal_out[497]) );
  DFFRHQX1 cal_out_reg_4__17_ ( .D(n1994), .CK(clk), .RN(rst_n), .Q(
        cal_out[417]) );
  DFFRHQX1 cal_out_reg_6__17_ ( .D(n2074), .CK(clk), .RN(rst_n), .Q(
        cal_out[337]) );
  DFFRHQX1 cal_out_reg_12__17_ ( .D(n2314), .CK(clk), .RN(rst_n), .Q(
        cal_out[97]) );
  DFFRHQX1 cal_out_reg_14__17_ ( .D(n2394), .CK(clk), .RN(rst_n), .Q(
        cal_out[17]) );
  DFFRHQX1 cal_out_reg_4__18_ ( .D(n1993), .CK(clk), .RN(rst_n), .Q(
        cal_out[418]) );
  DFFRHQX1 cal_out_reg_6__18_ ( .D(n2073), .CK(clk), .RN(rst_n), .Q(
        cal_out[338]) );
  DFFRHQX1 cal_out_reg_4__19_ ( .D(n1992), .CK(clk), .RN(rst_n), .Q(
        cal_out[419]) );
  DFFRHQX1 cal_out_reg_6__19_ ( .D(n2072), .CK(clk), .RN(rst_n), .Q(
        cal_out[339]) );
  DFFRHQX1 cal_out_reg_0__20_ ( .D(n1831), .CK(clk), .RN(rst_n), .Q(
        cal_out[580]) );
  DFFRHQX1 cal_out_reg_2__20_ ( .D(n1911), .CK(clk), .RN(rst_n), .Q(
        cal_out[500]) );
  DFFRHQX1 cal_out_reg_4__20_ ( .D(n1991), .CK(clk), .RN(rst_n), .Q(
        cal_out[420]) );
  DFFRHQX1 cal_out_reg_6__20_ ( .D(n2071), .CK(clk), .RN(rst_n), .Q(
        cal_out[340]) );
  DFFRHQX1 cal_out_reg_12__20_ ( .D(n2311), .CK(clk), .RN(rst_n), .Q(
        cal_out[100]) );
  DFFRHQX1 cal_out_reg_14__20_ ( .D(n2391), .CK(clk), .RN(rst_n), .Q(
        cal_out[20]) );
  DFFRHQX1 cal_out_reg_0__21_ ( .D(n1830), .CK(clk), .RN(rst_n), .Q(
        cal_out[581]) );
  DFFRHQX1 cal_out_reg_2__21_ ( .D(n1910), .CK(clk), .RN(rst_n), .Q(
        cal_out[501]) );
  DFFRHQX1 cal_out_reg_4__21_ ( .D(n1990), .CK(clk), .RN(rst_n), .Q(
        cal_out[421]) );
  DFFRHQX1 cal_out_reg_6__21_ ( .D(n2070), .CK(clk), .RN(rst_n), .Q(
        cal_out[341]) );
  DFFRHQX1 cal_out_reg_12__21_ ( .D(n2310), .CK(clk), .RN(rst_n), .Q(
        cal_out[101]) );
  DFFRHQX1 cal_out_reg_14__21_ ( .D(n2390), .CK(clk), .RN(rst_n), .Q(
        cal_out[21]) );
  DFFRHQX1 cal_out_reg_0__22_ ( .D(n1829), .CK(clk), .RN(rst_n), .Q(
        cal_out[582]) );
  DFFRHQX1 cal_out_reg_2__22_ ( .D(n1909), .CK(clk), .RN(rst_n), .Q(
        cal_out[502]) );
  DFFRHQX1 cal_out_reg_4__22_ ( .D(n1989), .CK(clk), .RN(rst_n), .Q(
        cal_out[422]) );
  DFFRHQX1 cal_out_reg_6__22_ ( .D(n2069), .CK(clk), .RN(rst_n), .Q(
        cal_out[342]) );
  DFFRHQX1 cal_out_reg_12__22_ ( .D(n2309), .CK(clk), .RN(rst_n), .Q(
        cal_out[102]) );
  DFFRHQX1 cal_out_reg_14__22_ ( .D(n2389), .CK(clk), .RN(rst_n), .Q(
        cal_out[22]) );
  DFFRHQX1 cal_out_reg_0__23_ ( .D(n1828), .CK(clk), .RN(rst_n), .Q(
        cal_out[583]) );
  DFFRHQX1 cal_out_reg_2__23_ ( .D(n1908), .CK(clk), .RN(rst_n), .Q(
        cal_out[503]) );
  DFFRHQX1 cal_out_reg_4__23_ ( .D(n1988), .CK(clk), .RN(rst_n), .Q(
        cal_out[423]) );
  DFFRHQX1 cal_out_reg_6__23_ ( .D(n2068), .CK(clk), .RN(rst_n), .Q(
        cal_out[343]) );
  DFFRHQX1 cal_out_reg_12__23_ ( .D(n2308), .CK(clk), .RN(rst_n), .Q(
        cal_out[103]) );
  DFFRHQX1 cal_out_reg_14__23_ ( .D(n2388), .CK(clk), .RN(rst_n), .Q(
        cal_out[23]) );
  DFFRHQX1 cal_out_reg_0__24_ ( .D(n1827), .CK(clk), .RN(rst_n), .Q(
        cal_out[584]) );
  DFFRHQX1 cal_out_reg_2__24_ ( .D(n1907), .CK(clk), .RN(rst_n), .Q(
        cal_out[504]) );
  DFFRHQX1 cal_out_reg_4__24_ ( .D(n1987), .CK(clk), .RN(rst_n), .Q(
        cal_out[424]) );
  DFFRHQX1 cal_out_reg_6__24_ ( .D(n2067), .CK(clk), .RN(rst_n), .Q(
        cal_out[344]) );
  DFFRHQX1 cal_out_reg_12__24_ ( .D(n2307), .CK(clk), .RN(rst_n), .Q(
        cal_out[104]) );
  DFFRHQX1 cal_out_reg_14__24_ ( .D(n2387), .CK(clk), .RN(rst_n), .Q(
        cal_out[24]) );
  DFFRHQX1 cal_out_reg_0__25_ ( .D(n1826), .CK(clk), .RN(rst_n), .Q(
        cal_out[585]) );
  DFFRHQX1 cal_out_reg_2__25_ ( .D(n1906), .CK(clk), .RN(rst_n), .Q(
        cal_out[505]) );
  DFFRHQX1 cal_out_reg_4__25_ ( .D(n1986), .CK(clk), .RN(rst_n), .Q(
        cal_out[425]) );
  DFFRHQX1 cal_out_reg_6__25_ ( .D(n2066), .CK(clk), .RN(rst_n), .Q(
        cal_out[345]) );
  DFFRHQX1 cal_out_reg_12__25_ ( .D(n2306), .CK(clk), .RN(rst_n), .Q(
        cal_out[105]) );
  DFFRHQX1 cal_out_reg_14__25_ ( .D(n2386), .CK(clk), .RN(rst_n), .Q(
        cal_out[25]) );
  DFFRHQX1 cal_out_reg_4__26_ ( .D(n1985), .CK(clk), .RN(rst_n), .Q(
        cal_out[426]) );
  DFFRHQX1 cal_out_reg_6__26_ ( .D(n2065), .CK(clk), .RN(rst_n), .Q(
        cal_out[346]) );
  DFFRHQX1 cal_out_reg_4__27_ ( .D(n1984), .CK(clk), .RN(rst_n), .Q(
        cal_out[427]) );
  DFFRHQX1 cal_out_reg_6__27_ ( .D(n2064), .CK(clk), .RN(rst_n), .Q(
        cal_out[347]) );
  DFFRHQX1 cal_out_reg_0__28_ ( .D(n1823), .CK(clk), .RN(rst_n), .Q(
        cal_out[588]) );
  DFFRHQX1 cal_out_reg_2__28_ ( .D(n1903), .CK(clk), .RN(rst_n), .Q(
        cal_out[508]) );
  DFFRHQX1 cal_out_reg_4__28_ ( .D(n1983), .CK(clk), .RN(rst_n), .Q(
        cal_out[428]) );
  DFFRHQX1 cal_out_reg_6__28_ ( .D(n2063), .CK(clk), .RN(rst_n), .Q(
        cal_out[348]) );
  DFFRHQX1 cal_out_reg_12__28_ ( .D(n2303), .CK(clk), .RN(rst_n), .Q(
        cal_out[108]) );
  DFFRHQX1 cal_out_reg_14__28_ ( .D(n2383), .CK(clk), .RN(rst_n), .Q(
        cal_out[28]) );
  DFFRHQX1 cal_out_reg_0__29_ ( .D(n1822), .CK(clk), .RN(rst_n), .Q(
        cal_out[589]) );
  DFFRHQX1 cal_out_reg_2__29_ ( .D(n1902), .CK(clk), .RN(rst_n), .Q(
        cal_out[509]) );
  DFFRHQX1 cal_out_reg_4__29_ ( .D(n1982), .CK(clk), .RN(rst_n), .Q(
        cal_out[429]) );
  DFFRHQX1 cal_out_reg_6__29_ ( .D(n2062), .CK(clk), .RN(rst_n), .Q(
        cal_out[349]) );
  DFFRHQX1 cal_out_reg_12__29_ ( .D(n2302), .CK(clk), .RN(rst_n), .Q(
        cal_out[109]) );
  DFFRHQX1 cal_out_reg_14__29_ ( .D(n2382), .CK(clk), .RN(rst_n), .Q(
        cal_out[29]) );
  DFFRHQX1 cal_out_reg_0__30_ ( .D(n1821), .CK(clk), .RN(rst_n), .Q(
        cal_out[590]) );
  DFFRHQX1 cal_out_reg_2__30_ ( .D(n1901), .CK(clk), .RN(rst_n), .Q(
        cal_out[510]) );
  DFFRHQX1 cal_out_reg_4__30_ ( .D(n1981), .CK(clk), .RN(rst_n), .Q(
        cal_out[430]) );
  DFFRHQX1 cal_out_reg_6__30_ ( .D(n2061), .CK(clk), .RN(rst_n), .Q(
        cal_out[350]) );
  DFFRHQX1 cal_out_reg_12__30_ ( .D(n2301), .CK(clk), .RN(rst_n), .Q(
        cal_out[110]) );
  DFFRHQX1 cal_out_reg_14__30_ ( .D(n2381), .CK(clk), .RN(rst_n), .Q(
        cal_out[30]) );
  DFFRHQX1 cal_out_reg_0__31_ ( .D(n1820), .CK(clk), .RN(rst_n), .Q(
        cal_out[591]) );
  DFFRHQX1 cal_out_reg_2__31_ ( .D(n1900), .CK(clk), .RN(rst_n), .Q(
        cal_out[511]) );
  DFFRHQX1 cal_out_reg_4__31_ ( .D(n1980), .CK(clk), .RN(rst_n), .Q(
        cal_out[431]) );
  DFFRHQX1 cal_out_reg_6__31_ ( .D(n2060), .CK(clk), .RN(rst_n), .Q(
        cal_out[351]) );
  DFFRHQX1 cal_out_reg_12__31_ ( .D(n2300), .CK(clk), .RN(rst_n), .Q(
        cal_out[111]) );
  DFFRHQX1 cal_out_reg_14__31_ ( .D(n2380), .CK(clk), .RN(rst_n), .Q(
        cal_out[31]) );
  DFFRHQX1 cal_out_reg_0__32_ ( .D(n1819), .CK(clk), .RN(rst_n), .Q(
        cal_out[592]) );
  DFFRHQX1 cal_out_reg_2__32_ ( .D(n1899), .CK(clk), .RN(rst_n), .Q(
        cal_out[512]) );
  DFFRHQX1 cal_out_reg_12__32_ ( .D(n2299), .CK(clk), .RN(rst_n), .Q(
        cal_out[112]) );
  DFFRHQX1 cal_out_reg_14__32_ ( .D(n2379), .CK(clk), .RN(rst_n), .Q(
        cal_out[32]) );
  DFFRHQX1 cal_out_reg_0__33_ ( .D(n1818), .CK(clk), .RN(rst_n), .Q(
        cal_out[593]) );
  DFFRHQX1 cal_out_reg_2__33_ ( .D(n1898), .CK(clk), .RN(rst_n), .Q(
        cal_out[513]) );
  DFFRHQX1 cal_out_reg_4__33_ ( .D(n1978), .CK(clk), .RN(rst_n), .Q(
        cal_out[433]) );
  DFFRHQX1 cal_out_reg_6__33_ ( .D(n2058), .CK(clk), .RN(rst_n), .Q(
        cal_out[353]) );
  DFFRHQX1 cal_out_reg_12__33_ ( .D(n2298), .CK(clk), .RN(rst_n), .Q(
        cal_out[113]) );
  DFFRHQX1 cal_out_reg_14__33_ ( .D(n2378), .CK(clk), .RN(rst_n), .Q(
        cal_out[33]) );
  DFFRHQX1 cal_out_reg_0__34_ ( .D(n1817), .CK(clk), .RN(rst_n), .Q(
        cal_out[594]) );
  DFFRHQX1 cal_out_reg_2__34_ ( .D(n1897), .CK(clk), .RN(rst_n), .Q(
        cal_out[514]) );
  DFFRHQX1 cal_out_reg_4__34_ ( .D(n1977), .CK(clk), .RN(rst_n), .Q(
        cal_out[434]) );
  DFFRHQX1 cal_out_reg_6__34_ ( .D(n2057), .CK(clk), .RN(rst_n), .Q(
        cal_out[354]) );
  DFFRHQX1 cal_out_reg_12__34_ ( .D(n2297), .CK(clk), .RN(rst_n), .Q(
        cal_out[114]) );
  DFFRHQX1 cal_out_reg_14__34_ ( .D(n2377), .CK(clk), .RN(rst_n), .Q(
        cal_out[34]) );
  DFFRHQX1 cal_out_reg_0__35_ ( .D(n1816), .CK(clk), .RN(rst_n), .Q(
        cal_out[595]) );
  DFFRHQX1 cal_out_reg_2__35_ ( .D(n1896), .CK(clk), .RN(rst_n), .Q(
        cal_out[515]) );
  DFFRHQX1 cal_out_reg_4__35_ ( .D(n1976), .CK(clk), .RN(rst_n), .Q(
        cal_out[435]) );
  DFFRHQX1 cal_out_reg_6__35_ ( .D(n2056), .CK(clk), .RN(rst_n), .Q(
        cal_out[355]) );
  DFFRHQX1 cal_out_reg_12__35_ ( .D(n2296), .CK(clk), .RN(rst_n), .Q(
        cal_out[115]) );
  DFFRHQX1 cal_out_reg_14__35_ ( .D(n2376), .CK(clk), .RN(rst_n), .Q(
        cal_out[35]) );
  DFFRHQX1 cal_out_reg_0__36_ ( .D(n1815), .CK(clk), .RN(rst_n), .Q(
        cal_out[596]) );
  DFFRHQX1 cal_out_reg_2__36_ ( .D(n1895), .CK(clk), .RN(rst_n), .Q(
        cal_out[516]) );
  DFFRHQX1 cal_out_reg_4__36_ ( .D(n1975), .CK(clk), .RN(rst_n), .Q(
        cal_out[436]) );
  DFFRHQX1 cal_out_reg_6__36_ ( .D(n2055), .CK(clk), .RN(rst_n), .Q(
        cal_out[356]) );
  DFFRHQX1 cal_out_reg_12__36_ ( .D(n2295), .CK(clk), .RN(rst_n), .Q(
        cal_out[116]) );
  DFFRHQX1 cal_out_reg_14__36_ ( .D(n2375), .CK(clk), .RN(rst_n), .Q(
        cal_out[36]) );
  DFFRHQX1 cal_out_reg_0__37_ ( .D(n1814), .CK(clk), .RN(rst_n), .Q(
        cal_out[597]) );
  DFFRHQX1 cal_out_reg_2__37_ ( .D(n1894), .CK(clk), .RN(rst_n), .Q(
        cal_out[517]) );
  DFFRHQX1 cal_out_reg_4__37_ ( .D(n1974), .CK(clk), .RN(rst_n), .Q(
        cal_out[437]) );
  DFFRHQX1 cal_out_reg_6__37_ ( .D(n2054), .CK(clk), .RN(rst_n), .Q(
        cal_out[357]) );
  DFFRHQX1 cal_out_reg_12__37_ ( .D(n2294), .CK(clk), .RN(rst_n), .Q(
        cal_out[117]) );
  DFFRHQX1 cal_out_reg_14__37_ ( .D(n2374), .CK(clk), .RN(rst_n), .Q(
        cal_out[37]) );
  DFFRHQX1 cal_out_reg_0__38_ ( .D(n1813), .CK(clk), .RN(rst_n), .Q(
        cal_out[598]) );
  DFFRHQX1 cal_out_reg_2__38_ ( .D(n1893), .CK(clk), .RN(rst_n), .Q(
        cal_out[518]) );
  DFFRHQX1 cal_out_reg_4__38_ ( .D(n1973), .CK(clk), .RN(rst_n), .Q(
        cal_out[438]) );
  DFFRHQX1 cal_out_reg_6__38_ ( .D(n2053), .CK(clk), .RN(rst_n), .Q(
        cal_out[358]) );
  DFFRHQX1 cal_out_reg_12__38_ ( .D(n2293), .CK(clk), .RN(rst_n), .Q(
        cal_out[118]) );
  DFFRHQX1 cal_out_reg_14__38_ ( .D(n2373), .CK(clk), .RN(rst_n), .Q(
        cal_out[38]) );
  DFFRHQX1 cal_out_reg_0__39_ ( .D(n1812), .CK(clk), .RN(rst_n), .Q(
        cal_out[599]) );
  DFFRHQX1 cal_out_reg_2__39_ ( .D(n1892), .CK(clk), .RN(rst_n), .Q(
        cal_out[519]) );
  DFFRHQX1 cal_out_reg_4__39_ ( .D(n1972), .CK(clk), .RN(rst_n), .Q(
        cal_out[439]) );
  DFFRHQX1 cal_out_reg_6__39_ ( .D(n2052), .CK(clk), .RN(rst_n), .Q(
        cal_out[359]) );
  DFFRHQX1 cal_out_reg_12__39_ ( .D(n2292), .CK(clk), .RN(rst_n), .Q(
        cal_out[119]) );
  DFFRHQX1 cal_out_reg_14__39_ ( .D(n2372), .CK(clk), .RN(rst_n), .Q(
        cal_out[39]) );
  DFFRHQX1 length_reg_reg_0__5_ ( .D(n1722), .CK(clk), .RN(rst_n), .Q(
        length_reg[89]) );
  DFFRHQX1 length_reg_reg_2__5_ ( .D(n1734), .CK(clk), .RN(rst_n), .Q(
        length_reg[77]) );
  DFFRHQX1 length_reg_reg_12__5_ ( .D(n1794), .CK(clk), .RN(rst_n), .Q(
        length_reg[17]) );
  DFFRHQX1 length_reg_reg_14__5_ ( .D(n1806), .CK(clk), .RN(rst_n), .Q(
        length_reg[5]) );
  DFFRHQX1 length_reg_reg_0__3_ ( .D(n1724), .CK(clk), .RN(rst_n), .Q(
        length_reg[87]) );
  DFFRHQX1 length_reg_reg_2__3_ ( .D(n1736), .CK(clk), .RN(rst_n), .Q(
        length_reg[75]) );
  DFFRHQX1 length_reg_reg_4__3_ ( .D(n1748), .CK(clk), .RN(rst_n), .Q(
        length_reg[63]) );
  DFFRHQX1 length_reg_reg_6__3_ ( .D(n1760), .CK(clk), .RN(rst_n), .Q(
        length_reg[51]) );
  DFFRHQX1 length_reg_reg_12__3_ ( .D(n1796), .CK(clk), .RN(rst_n), .Q(
        length_reg[15]) );
  DFFRHQX1 length_reg_reg_14__3_ ( .D(n1808), .CK(clk), .RN(rst_n), .Q(
        length_reg[3]) );
  DFFRHQX1 length_reg_reg_0__1_ ( .D(n1726), .CK(clk), .RN(rst_n), .Q(
        length_reg[85]) );
  DFFRHQX1 length_reg_reg_2__1_ ( .D(n1738), .CK(clk), .RN(rst_n), .Q(
        length_reg[73]) );
  DFFRHQX1 length_reg_reg_4__1_ ( .D(n1750), .CK(clk), .RN(rst_n), .Q(
        length_reg[61]) );
  DFFRHQX1 length_reg_reg_6__1_ ( .D(n1762), .CK(clk), .RN(rst_n), .Q(
        length_reg[49]) );
  DFFRHQX1 length_reg_reg_12__1_ ( .D(n1798), .CK(clk), .RN(rst_n), .Q(
        length_reg[13]) );
  DFFRHQX1 length_reg_reg_14__1_ ( .D(n1810), .CK(clk), .RN(rst_n), .Q(
        length_reg[1]) );
  DFFRHQX1 length_reg_reg_0__4_ ( .D(n1723), .CK(clk), .RN(rst_n), .Q(
        length_reg[88]) );
  DFFRHQX1 length_reg_reg_2__4_ ( .D(n1735), .CK(clk), .RN(rst_n), .Q(
        length_reg[76]) );
  DFFRHQX1 length_reg_reg_4__4_ ( .D(n1747), .CK(clk), .RN(rst_n), .Q(
        length_reg[64]) );
  DFFRHQX1 length_reg_reg_6__4_ ( .D(n1759), .CK(clk), .RN(rst_n), .Q(
        length_reg[52]) );
  DFFRHQX1 length_reg_reg_12__4_ ( .D(n1795), .CK(clk), .RN(rst_n), .Q(
        length_reg[16]) );
  DFFRHQX1 length_reg_reg_14__4_ ( .D(n1807), .CK(clk), .RN(rst_n), .Q(
        length_reg[4]) );
  DFFRHQX1 length_reg_reg_0__2_ ( .D(n1725), .CK(clk), .RN(rst_n), .Q(
        length_reg[86]) );
  DFFRHQX1 length_reg_reg_2__2_ ( .D(n1737), .CK(clk), .RN(rst_n), .Q(
        length_reg[74]) );
  DFFRHQX1 length_reg_reg_4__2_ ( .D(n1749), .CK(clk), .RN(rst_n), .Q(
        length_reg[62]) );
  DFFRHQX1 length_reg_reg_6__2_ ( .D(n1761), .CK(clk), .RN(rst_n), .Q(
        length_reg[50]) );
  DFFRHQX1 length_reg_reg_12__2_ ( .D(n1797), .CK(clk), .RN(rst_n), .Q(
        length_reg[14]) );
  DFFRHQX1 length_reg_reg_14__2_ ( .D(n1809), .CK(clk), .RN(rst_n), .Q(
        length_reg[2]) );
  DFFRHQX1 length_reg_reg_0__0_ ( .D(n1727), .CK(clk), .RN(rst_n), .Q(
        length_reg[84]) );
  DFFRHQX1 length_reg_reg_2__0_ ( .D(n1739), .CK(clk), .RN(rst_n), .Q(
        length_reg[72]) );
  DFFRHQX1 length_reg_reg_4__0_ ( .D(n1751), .CK(clk), .RN(rst_n), .Q(
        length_reg[60]) );
  DFFRHQX1 length_reg_reg_6__0_ ( .D(n1763), .CK(clk), .RN(rst_n), .Q(
        length_reg[48]) );
  DFFRHQX1 length_reg_reg_12__0_ ( .D(n1799), .CK(clk), .RN(rst_n), .Q(
        length_reg[12]) );
  DFFRHQX1 length_reg_reg_14__0_ ( .D(n1811), .CK(clk), .RN(rst_n), .Q(
        length_reg[0]) );
  DFFRHQX1 cal_out_reg_10__0_ ( .D(n2251), .CK(clk), .RN(rst_n), .Q(
        cal_out[160]) );
  DFFRHQX1 cal_out_reg_10__1_ ( .D(n2250), .CK(clk), .RN(rst_n), .Q(
        cal_out[161]) );
  DFFRHQX1 cal_out_reg_10__4_ ( .D(n2247), .CK(clk), .RN(rst_n), .Q(
        cal_out[164]) );
  DFFRHQX1 cal_out_reg_10__5_ ( .D(n2246), .CK(clk), .RN(rst_n), .Q(
        cal_out[165]) );
  DFFRHQX1 cal_out_reg_10__6_ ( .D(n2245), .CK(clk), .RN(rst_n), .Q(
        cal_out[166]) );
  DFFRHQX1 cal_out_reg_10__7_ ( .D(n2244), .CK(clk), .RN(rst_n), .Q(
        cal_out[167]) );
  DFFRHQX1 cal_out_reg_10__8_ ( .D(n2243), .CK(clk), .RN(rst_n), .Q(
        cal_out[168]) );
  DFFRHQX1 cal_out_reg_10__9_ ( .D(n2242), .CK(clk), .RN(rst_n), .Q(
        cal_out[169]) );
  DFFRHQX1 cal_out_reg_10__12_ ( .D(n2239), .CK(clk), .RN(rst_n), .Q(
        cal_out[172]) );
  DFFRHQX1 cal_out_reg_10__13_ ( .D(n2238), .CK(clk), .RN(rst_n), .Q(
        cal_out[173]) );
  DFFRHQX1 cal_out_reg_10__14_ ( .D(n2237), .CK(clk), .RN(rst_n), .Q(
        cal_out[174]) );
  DFFRHQX1 cal_out_reg_10__15_ ( .D(n2236), .CK(clk), .RN(rst_n), .Q(
        cal_out[175]) );
  DFFRHQX1 cal_out_reg_10__16_ ( .D(n2235), .CK(clk), .RN(rst_n), .Q(
        cal_out[176]) );
  DFFRHQX1 cal_out_reg_10__17_ ( .D(n2234), .CK(clk), .RN(rst_n), .Q(
        cal_out[177]) );
  DFFRHQX1 cal_out_reg_10__18_ ( .D(n2233), .CK(clk), .RN(rst_n), .Q(
        cal_out[178]) );
  DFFRHQX1 cal_out_reg_10__19_ ( .D(n2232), .CK(clk), .RN(rst_n), .Q(
        cal_out[179]) );
  DFFRHQX1 cal_out_reg_10__20_ ( .D(n2231), .CK(clk), .RN(rst_n), .Q(
        cal_out[180]) );
  DFFRHQX1 cal_out_reg_10__21_ ( .D(n2230), .CK(clk), .RN(rst_n), .Q(
        cal_out[181]) );
  DFFRHQX1 cal_out_reg_10__22_ ( .D(n2229), .CK(clk), .RN(rst_n), .Q(
        cal_out[182]) );
  DFFRHQX1 cal_out_reg_10__23_ ( .D(n2228), .CK(clk), .RN(rst_n), .Q(
        cal_out[183]) );
  DFFRHQX1 cal_out_reg_10__24_ ( .D(n2227), .CK(clk), .RN(rst_n), .Q(
        cal_out[184]) );
  DFFRHQX1 cal_out_reg_10__25_ ( .D(n2226), .CK(clk), .RN(rst_n), .Q(
        cal_out[185]) );
  DFFRHQX1 cal_out_reg_10__26_ ( .D(n2225), .CK(clk), .RN(rst_n), .Q(
        cal_out[186]) );
  DFFRHQX1 cal_out_reg_10__27_ ( .D(n2224), .CK(clk), .RN(rst_n), .Q(
        cal_out[187]) );
  DFFRHQX1 cal_out_reg_10__28_ ( .D(n2223), .CK(clk), .RN(rst_n), .Q(
        cal_out[188]) );
  DFFRHQX1 cal_out_reg_10__29_ ( .D(n2222), .CK(clk), .RN(rst_n), .Q(
        cal_out[189]) );
  DFFRHQX1 cal_out_reg_10__30_ ( .D(n2221), .CK(clk), .RN(rst_n), .Q(
        cal_out[190]) );
  DFFRHQX1 cal_out_reg_10__31_ ( .D(n2220), .CK(clk), .RN(rst_n), .Q(
        cal_out[191]) );
  DFFRHQX1 cal_out_reg_10__33_ ( .D(n2218), .CK(clk), .RN(rst_n), .Q(
        cal_out[193]) );
  DFFRHQX1 cal_out_reg_10__34_ ( .D(n2217), .CK(clk), .RN(rst_n), .Q(
        cal_out[194]) );
  DFFRHQX1 cal_out_reg_10__35_ ( .D(n2216), .CK(clk), .RN(rst_n), .Q(
        cal_out[195]) );
  DFFRHQX1 cal_out_reg_10__36_ ( .D(n2215), .CK(clk), .RN(rst_n), .Q(
        cal_out[196]) );
  DFFRHQX1 cal_out_reg_10__37_ ( .D(n2214), .CK(clk), .RN(rst_n), .Q(
        cal_out[197]) );
  DFFRHQX1 cal_out_reg_10__38_ ( .D(n2213), .CK(clk), .RN(rst_n), .Q(
        cal_out[198]) );
  DFFRHQX1 cal_out_reg_10__39_ ( .D(n2212), .CK(clk), .RN(rst_n), .Q(
        cal_out[199]) );
  DFFRHQX1 length_reg_reg_10__5_ ( .D(n1782), .CK(clk), .RN(rst_n), .Q(
        length_reg[29]) );
  DFFRHQX1 length_reg_reg_10__3_ ( .D(n1784), .CK(clk), .RN(rst_n), .Q(
        length_reg[27]) );
  DFFRHQX1 length_reg_reg_10__1_ ( .D(n1786), .CK(clk), .RN(rst_n), .Q(
        length_reg[25]) );
  DFFRHQX1 length_reg_reg_10__4_ ( .D(n1783), .CK(clk), .RN(rst_n), .Q(
        length_reg[28]) );
  DFFRHQX1 length_reg_reg_10__2_ ( .D(n1785), .CK(clk), .RN(rst_n), .Q(
        length_reg[26]) );
  DFFRHQX1 length_reg_reg_10__0_ ( .D(n1787), .CK(clk), .RN(rst_n), .Q(
        length_reg[24]) );
  DFFRHQX1 i_mat_reg_3_ ( .D(N1289), .CK(clk), .RN(rst_n), .Q(i_mat[3]) );
  DFFRHQX1 w_mat_reg_3_ ( .D(N1294), .CK(clk), .RN(rst_n), .Q(w_mat[3]) );
  DFFRHQX1 cal_cnt_reg_7_ ( .D(N11321), .CK(clk), .RN(rst_n), .Q(cal_cnt[7])
         );
  DFFRHQX1 i_mat_reg_0_ ( .D(N1286), .CK(clk), .RN(rst_n), .Q(i_mat[0]) );
  DFFRHQX1 i_mat_reg_1_ ( .D(N1287), .CK(clk), .RN(rst_n), .Q(i_mat[1]) );
  DFFRHQX1 i_mat_reg_2_ ( .D(N1288), .CK(clk), .RN(rst_n), .Q(i_mat[2]) );
  DFFRHQX1 w_mat_reg_0_ ( .D(N1291), .CK(clk), .RN(rst_n), .Q(w_mat[0]) );
  DFFRHQX1 w_mat_reg_1_ ( .D(N1292), .CK(clk), .RN(rst_n), .Q(w_mat[1]) );
  DFFRHQX1 w_mat_reg_2_ ( .D(N1293), .CK(clk), .RN(rst_n), .Q(w_mat[2]) );
  DFFRHQX1 cal_cnt_reg_3_ ( .D(N11317), .CK(clk), .RN(rst_n), .Q(cal_cnt[3])
         );
  DFFRHQX1 c_plus_reg_14_ ( .D(N12580), .CK(clk), .RN(rst_n), .Q(c_plus[14])
         );
  DFFRHQX1 in_cnt_reg_7_ ( .D(n5824), .CK(clk), .RN(rst_n), .Q(in_cnt[7]) );
  DFFRHQX1 c_plus_reg_30_ ( .D(N12596), .CK(clk), .RN(rst_n), .Q(c_plus[30])
         );
  DFFRHQX1 in_cnt_64_reg_5_ ( .D(N1045), .CK(clk), .RN(rst_n), .Q(in_cnt_64[5]) );
  DFFRHQX1 c_plus_reg_6_ ( .D(N12572), .CK(clk), .RN(rst_n), .Q(c_plus[6]) );
  DFFRHQX1 c_plus_reg_3_ ( .D(N12569), .CK(clk), .RN(rst_n), .Q(c_plus[3]) );
  DFFRHQX1 cal_out_reg_1__1_ ( .D(n1890), .CK(clk), .RN(rst_n), .Q(
        cal_out[521]) );
  DFFRHQX1 cal_out_reg_3__1_ ( .D(n1970), .CK(clk), .RN(rst_n), .Q(
        cal_out[441]) );
  DFFRHQX1 cal_out_reg_7__1_ ( .D(n2130), .CK(clk), .RN(rst_n), .Q(
        cal_out[281]) );
  DFFRHQX1 cal_out_reg_13__1_ ( .D(n2370), .CK(clk), .RN(rst_n), .Q(
        cal_out[41]) );
  DFFRHQX1 cal_out_reg_1__2_ ( .D(n1889), .CK(clk), .RN(rst_n), .Q(
        cal_out[522]) );
  DFFRHQX1 cal_out_reg_3__2_ ( .D(n1969), .CK(clk), .RN(rst_n), .Q(
        cal_out[442]) );
  DFFRHQX1 cal_out_reg_5__2_ ( .D(n2049), .CK(clk), .RN(rst_n), .Q(
        cal_out[362]) );
  DFFRHQX1 cal_out_reg_7__2_ ( .D(n2129), .CK(clk), .RN(rst_n), .Q(
        cal_out[282]) );
  DFFRHQX1 cal_out_reg_11__2_ ( .D(n2289), .CK(clk), .RN(rst_n), .Q(
        cal_out[122]) );
  DFFRHQX1 cal_out_reg_13__2_ ( .D(n2369), .CK(clk), .RN(rst_n), .Q(
        cal_out[42]) );
  DFFRHQX1 cal_out_reg_1__3_ ( .D(n1888), .CK(clk), .RN(rst_n), .Q(
        cal_out[523]) );
  DFFRHQX1 cal_out_reg_3__3_ ( .D(n1968), .CK(clk), .RN(rst_n), .Q(
        cal_out[443]) );
  DFFRHQX1 cal_out_reg_7__3_ ( .D(n2128), .CK(clk), .RN(rst_n), .Q(
        cal_out[283]) );
  DFFRHQX1 cal_out_reg_13__3_ ( .D(n2368), .CK(clk), .RN(rst_n), .Q(
        cal_out[43]) );
  DFFRHQX1 cal_out_reg_1__5_ ( .D(n1886), .CK(clk), .RN(rst_n), .Q(
        cal_out[525]) );
  DFFRHQX1 cal_out_reg_3__5_ ( .D(n1966), .CK(clk), .RN(rst_n), .Q(
        cal_out[445]) );
  DFFRHQX1 cal_out_reg_7__5_ ( .D(n2126), .CK(clk), .RN(rst_n), .Q(
        cal_out[285]) );
  DFFRHQX1 cal_out_reg_13__5_ ( .D(n2366), .CK(clk), .RN(rst_n), .Q(
        cal_out[45]) );
  DFFRHQX1 cal_out_reg_1__7_ ( .D(n1884), .CK(clk), .RN(rst_n), .Q(
        cal_out[527]) );
  DFFRHQX1 cal_out_reg_3__7_ ( .D(n1964), .CK(clk), .RN(rst_n), .Q(
        cal_out[447]) );
  DFFRHQX1 cal_out_reg_7__7_ ( .D(n2124), .CK(clk), .RN(rst_n), .Q(
        cal_out[287]) );
  DFFRHQX1 cal_out_reg_13__7_ ( .D(n2364), .CK(clk), .RN(rst_n), .Q(
        cal_out[47]) );
  DFFRHQX1 cal_out_reg_1__9_ ( .D(n1882), .CK(clk), .RN(rst_n), .Q(
        cal_out[529]) );
  DFFRHQX1 cal_out_reg_3__9_ ( .D(n1962), .CK(clk), .RN(rst_n), .Q(
        cal_out[449]) );
  DFFRHQX1 cal_out_reg_7__9_ ( .D(n2122), .CK(clk), .RN(rst_n), .Q(
        cal_out[289]) );
  DFFRHQX1 cal_out_reg_13__9_ ( .D(n2362), .CK(clk), .RN(rst_n), .Q(
        cal_out[49]) );
  DFFRHQX1 cal_out_reg_1__10_ ( .D(n1881), .CK(clk), .RN(rst_n), .Q(
        cal_out[530]) );
  DFFRHQX1 cal_out_reg_3__10_ ( .D(n1961), .CK(clk), .RN(rst_n), .Q(
        cal_out[450]) );
  DFFRHQX1 cal_out_reg_5__10_ ( .D(n2041), .CK(clk), .RN(rst_n), .Q(
        cal_out[370]) );
  DFFRHQX1 cal_out_reg_7__10_ ( .D(n2121), .CK(clk), .RN(rst_n), .Q(
        cal_out[290]) );
  DFFRHQX1 cal_out_reg_11__10_ ( .D(n2281), .CK(clk), .RN(rst_n), .Q(
        cal_out[130]) );
  DFFRHQX1 cal_out_reg_13__10_ ( .D(n2361), .CK(clk), .RN(rst_n), .Q(
        cal_out[50]) );
  DFFRHQX1 cal_out_reg_1__11_ ( .D(n1880), .CK(clk), .RN(rst_n), .Q(
        cal_out[531]) );
  DFFRHQX1 cal_out_reg_3__11_ ( .D(n1960), .CK(clk), .RN(rst_n), .Q(
        cal_out[451]) );
  DFFRHQX1 cal_out_reg_7__11_ ( .D(n2120), .CK(clk), .RN(rst_n), .Q(
        cal_out[291]) );
  DFFRHQX1 cal_out_reg_13__11_ ( .D(n2360), .CK(clk), .RN(rst_n), .Q(
        cal_out[51]) );
  DFFRHQX1 cal_out_reg_1__13_ ( .D(n1878), .CK(clk), .RN(rst_n), .Q(
        cal_out[533]) );
  DFFRHQX1 cal_out_reg_3__13_ ( .D(n1958), .CK(clk), .RN(rst_n), .Q(
        cal_out[453]) );
  DFFRHQX1 cal_out_reg_13__13_ ( .D(n2358), .CK(clk), .RN(rst_n), .Q(
        cal_out[53]) );
  DFFRHQX1 cal_out_reg_1__15_ ( .D(n1876), .CK(clk), .RN(rst_n), .Q(
        cal_out[535]) );
  DFFRHQX1 cal_out_reg_3__15_ ( .D(n1956), .CK(clk), .RN(rst_n), .Q(
        cal_out[455]) );
  DFFRHQX1 cal_out_reg_13__15_ ( .D(n2356), .CK(clk), .RN(rst_n), .Q(
        cal_out[55]) );
  DFFRHQX1 cal_out_reg_1__18_ ( .D(n1873), .CK(clk), .RN(rst_n), .Q(
        cal_out[538]) );
  DFFRHQX1 cal_out_reg_3__18_ ( .D(n1953), .CK(clk), .RN(rst_n), .Q(
        cal_out[458]) );
  DFFRHQX1 cal_out_reg_7__18_ ( .D(n2113), .CK(clk), .RN(rst_n), .Q(
        cal_out[298]) );
  DFFRHQX1 cal_out_reg_13__18_ ( .D(n2353), .CK(clk), .RN(rst_n), .Q(
        cal_out[58]) );
  DFFRHQX1 cal_out_reg_1__19_ ( .D(n1872), .CK(clk), .RN(rst_n), .Q(
        cal_out[539]) );
  DFFRHQX1 cal_out_reg_3__19_ ( .D(n1952), .CK(clk), .RN(rst_n), .Q(
        cal_out[459]) );
  DFFRHQX1 cal_out_reg_7__19_ ( .D(n2112), .CK(clk), .RN(rst_n), .Q(
        cal_out[299]) );
  DFFRHQX1 cal_out_reg_13__19_ ( .D(n2352), .CK(clk), .RN(rst_n), .Q(
        cal_out[59]) );
  DFFRHQX1 cal_out_reg_1__26_ ( .D(n1865), .CK(clk), .RN(rst_n), .Q(
        cal_out[546]) );
  DFFRHQX1 cal_out_reg_3__26_ ( .D(n1945), .CK(clk), .RN(rst_n), .Q(
        cal_out[466]) );
  DFFRHQX1 cal_out_reg_7__26_ ( .D(n2105), .CK(clk), .RN(rst_n), .Q(
        cal_out[306]) );
  DFFRHQX1 cal_out_reg_13__26_ ( .D(n2345), .CK(clk), .RN(rst_n), .Q(
        cal_out[66]) );
  DFFRHQX1 cal_out_reg_1__27_ ( .D(n1864), .CK(clk), .RN(rst_n), .Q(
        cal_out[547]) );
  DFFRHQX1 cal_out_reg_3__27_ ( .D(n1944), .CK(clk), .RN(rst_n), .Q(
        cal_out[467]) );
  DFFRHQX1 cal_out_reg_7__27_ ( .D(n2104), .CK(clk), .RN(rst_n), .Q(
        cal_out[307]) );
  DFFRHQX1 cal_out_reg_13__27_ ( .D(n2344), .CK(clk), .RN(rst_n), .Q(
        cal_out[67]) );
  DFFRHQX1 length_reg_reg_3__0_ ( .D(n1745), .CK(clk), .RN(rst_n), .Q(
        length_reg[66]) );
  DFFRHQX1 length_reg_reg_13__0_ ( .D(n1805), .CK(clk), .RN(rst_n), .Q(
        length_reg[6]) );
  DFFRHQX1 cal_out_reg_9__1_ ( .D(n2210), .CK(clk), .RN(rst_n), .Q(
        cal_out[201]) );
  DFFRHQX1 cal_out_reg_9__2_ ( .D(n2209), .CK(clk), .RN(rst_n), .Q(
        cal_out[202]) );
  DFFRHQX1 cal_out_reg_9__3_ ( .D(n2208), .CK(clk), .RN(rst_n), .Q(
        cal_out[203]) );
  DFFRHQX1 cal_out_reg_9__9_ ( .D(n2202), .CK(clk), .RN(rst_n), .Q(
        cal_out[209]) );
  DFFRHQX1 cal_out_reg_9__10_ ( .D(n2201), .CK(clk), .RN(rst_n), .Q(
        cal_out[210]) );
  DFFRHQX1 cal_out_reg_9__11_ ( .D(n2200), .CK(clk), .RN(rst_n), .Q(
        cal_out[211]) );
  DFFRHQX1 cal_out_reg_9__18_ ( .D(n2193), .CK(clk), .RN(rst_n), .Q(
        cal_out[218]) );
  DFFRHQX1 cal_out_reg_9__19_ ( .D(n2192), .CK(clk), .RN(rst_n), .Q(
        cal_out[219]) );
  DFFRHQX1 cal_out_reg_9__26_ ( .D(n2185), .CK(clk), .RN(rst_n), .Q(
        cal_out[226]) );
  DFFRHQX1 cal_out_reg_9__27_ ( .D(n2184), .CK(clk), .RN(rst_n), .Q(
        cal_out[227]) );
  DFFRHQX1 cal_out_reg_8__2_ ( .D(n2169), .CK(clk), .RN(rst_n), .Q(
        cal_out[242]) );
  DFFRHQX1 cal_out_reg_8__3_ ( .D(n2168), .CK(clk), .RN(rst_n), .Q(
        cal_out[243]) );
  DFFRHQX1 cal_out_reg_8__10_ ( .D(n2161), .CK(clk), .RN(rst_n), .Q(
        cal_out[250]) );
  DFFRHQX1 cal_out_reg_8__11_ ( .D(n2160), .CK(clk), .RN(rst_n), .Q(
        cal_out[251]) );
  DFFRHQX1 cal_out_reg_8__18_ ( .D(n2153), .CK(clk), .RN(rst_n), .Q(
        cal_out[258]) );
  DFFRHQX1 cal_out_reg_8__19_ ( .D(n2152), .CK(clk), .RN(rst_n), .Q(
        cal_out[259]) );
  DFFRHQX1 cal_out_reg_8__26_ ( .D(n2145), .CK(clk), .RN(rst_n), .Q(
        cal_out[266]) );
  DFFRHQX1 cal_out_reg_8__27_ ( .D(n2144), .CK(clk), .RN(rst_n), .Q(
        cal_out[267]) );
  DFFRHQX1 cal_out_reg_0__1_ ( .D(n1850), .CK(clk), .RN(rst_n), .Q(
        cal_out[561]) );
  DFFRHQX1 cal_out_reg_12__1_ ( .D(n2330), .CK(clk), .RN(rst_n), .Q(
        cal_out[81]) );
  DFFRHQX1 cal_out_reg_14__1_ ( .D(n2410), .CK(clk), .RN(rst_n), .Q(cal_out[1]) );
  DFFRHQX1 cal_out_reg_0__2_ ( .D(n1849), .CK(clk), .RN(rst_n), .Q(
        cal_out[562]) );
  DFFRHQX1 cal_out_reg_2__2_ ( .D(n1929), .CK(clk), .RN(rst_n), .Q(
        cal_out[482]) );
  DFFRHQX1 cal_out_reg_12__2_ ( .D(n2329), .CK(clk), .RN(rst_n), .Q(
        cal_out[82]) );
  DFFRHQX1 cal_out_reg_14__2_ ( .D(n2409), .CK(clk), .RN(rst_n), .Q(cal_out[2]) );
  DFFRHQX1 cal_out_reg_0__3_ ( .D(n1848), .CK(clk), .RN(rst_n), .Q(
        cal_out[563]) );
  DFFRHQX1 cal_out_reg_2__3_ ( .D(n1928), .CK(clk), .RN(rst_n), .Q(
        cal_out[483]) );
  DFFRHQX1 cal_out_reg_12__3_ ( .D(n2328), .CK(clk), .RN(rst_n), .Q(
        cal_out[83]) );
  DFFRHQX1 cal_out_reg_14__3_ ( .D(n2408), .CK(clk), .RN(rst_n), .Q(cal_out[3]) );
  DFFRHQX1 cal_out_reg_12__9_ ( .D(n2322), .CK(clk), .RN(rst_n), .Q(
        cal_out[89]) );
  DFFRHQX1 cal_out_reg_14__9_ ( .D(n2402), .CK(clk), .RN(rst_n), .Q(cal_out[9]) );
  DFFRHQX1 cal_out_reg_0__10_ ( .D(n1841), .CK(clk), .RN(rst_n), .Q(
        cal_out[570]) );
  DFFRHQX1 cal_out_reg_2__10_ ( .D(n1921), .CK(clk), .RN(rst_n), .Q(
        cal_out[490]) );
  DFFRHQX1 cal_out_reg_12__10_ ( .D(n2321), .CK(clk), .RN(rst_n), .Q(
        cal_out[90]) );
  DFFRHQX1 cal_out_reg_14__10_ ( .D(n2401), .CK(clk), .RN(rst_n), .Q(
        cal_out[10]) );
  DFFRHQX1 cal_out_reg_0__11_ ( .D(n1840), .CK(clk), .RN(rst_n), .Q(
        cal_out[571]) );
  DFFRHQX1 cal_out_reg_2__11_ ( .D(n1920), .CK(clk), .RN(rst_n), .Q(
        cal_out[491]) );
  DFFRHQX1 cal_out_reg_12__11_ ( .D(n2320), .CK(clk), .RN(rst_n), .Q(
        cal_out[91]) );
  DFFRHQX1 cal_out_reg_14__11_ ( .D(n2400), .CK(clk), .RN(rst_n), .Q(
        cal_out[11]) );
  DFFRHQX1 cal_out_reg_0__18_ ( .D(n1833), .CK(clk), .RN(rst_n), .Q(
        cal_out[578]) );
  DFFRHQX1 cal_out_reg_2__18_ ( .D(n1913), .CK(clk), .RN(rst_n), .Q(
        cal_out[498]) );
  DFFRHQX1 cal_out_reg_12__18_ ( .D(n2313), .CK(clk), .RN(rst_n), .Q(
        cal_out[98]) );
  DFFRHQX1 cal_out_reg_14__18_ ( .D(n2393), .CK(clk), .RN(rst_n), .Q(
        cal_out[18]) );
  DFFRHQX1 cal_out_reg_0__19_ ( .D(n1832), .CK(clk), .RN(rst_n), .Q(
        cal_out[579]) );
  DFFRHQX1 cal_out_reg_2__19_ ( .D(n1912), .CK(clk), .RN(rst_n), .Q(
        cal_out[499]) );
  DFFRHQX1 cal_out_reg_12__19_ ( .D(n2312), .CK(clk), .RN(rst_n), .Q(
        cal_out[99]) );
  DFFRHQX1 cal_out_reg_14__19_ ( .D(n2392), .CK(clk), .RN(rst_n), .Q(
        cal_out[19]) );
  DFFRHQX1 cal_out_reg_0__26_ ( .D(n1825), .CK(clk), .RN(rst_n), .Q(
        cal_out[586]) );
  DFFRHQX1 cal_out_reg_2__26_ ( .D(n1905), .CK(clk), .RN(rst_n), .Q(
        cal_out[506]) );
  DFFRHQX1 cal_out_reg_12__26_ ( .D(n2305), .CK(clk), .RN(rst_n), .Q(
        cal_out[106]) );
  DFFRHQX1 cal_out_reg_14__26_ ( .D(n2385), .CK(clk), .RN(rst_n), .Q(
        cal_out[26]) );
  DFFRHQX1 cal_out_reg_0__27_ ( .D(n1824), .CK(clk), .RN(rst_n), .Q(
        cal_out[587]) );
  DFFRHQX1 cal_out_reg_2__27_ ( .D(n1904), .CK(clk), .RN(rst_n), .Q(
        cal_out[507]) );
  DFFRHQX1 cal_out_reg_12__27_ ( .D(n2304), .CK(clk), .RN(rst_n), .Q(
        cal_out[107]) );
  DFFRHQX1 cal_out_reg_14__27_ ( .D(n2384), .CK(clk), .RN(rst_n), .Q(
        cal_out[27]) );
  DFFRHQX1 cal_out_reg_10__2_ ( .D(n2249), .CK(clk), .RN(rst_n), .Q(
        cal_out[162]) );
  DFFRHQX1 cal_out_reg_10__3_ ( .D(n2248), .CK(clk), .RN(rst_n), .Q(
        cal_out[163]) );
  DFFRHQX1 cal_out_reg_10__10_ ( .D(n2241), .CK(clk), .RN(rst_n), .Q(
        cal_out[170]) );
  DFFRHQX1 cal_out_reg_10__11_ ( .D(n2240), .CK(clk), .RN(rst_n), .Q(
        cal_out[171]) );
  DFFRHQX1 calin_cnt_reg_7_ ( .D(N1369), .CK(clk), .RN(rst_n), .Q(calin_cnt[7]) );
  DFFRHQX1 cal_cnt_reg_1_ ( .D(N11315), .CK(clk), .RN(rst_n), .Q(cal_cnt[1])
         );
  DFFRHQX1 cal_cnt_reg_2_ ( .D(N11316), .CK(clk), .RN(rst_n), .Q(cal_cnt[2])
         );
  DFFRHQX1 out_cnt_reg_5_ ( .D(n5834), .CK(clk), .RN(rst_n), .Q(out_cnt[5]) );
  DFFRHQX1 c_plus_reg_11_ ( .D(N12577), .CK(clk), .RN(rst_n), .Q(c_plus[11])
         );
  DFFRHQX1 c_plus_reg_12_ ( .D(N12578), .CK(clk), .RN(rst_n), .Q(c_plus[12])
         );
  DFFRHQX1 c_plus_reg_8_ ( .D(N12574), .CK(clk), .RN(rst_n), .Q(c_plus[8]) );
  DFFRHQX1 c_plus_reg_10_ ( .D(N12576), .CK(clk), .RN(rst_n), .Q(c_plus[10])
         );
  DFFRHQX1 c_plus_reg_9_ ( .D(N12575), .CK(clk), .RN(rst_n), .Q(c_plus[9]) );
  DFFRHQX1 c_plus_reg_7_ ( .D(N12573), .CK(clk), .RN(rst_n), .Q(c_plus[7]) );
  DFFRHQX1 out_cnt_reg_4_ ( .D(n5835), .CK(clk), .RN(rst_n), .Q(out_cnt[4]) );
  DFFRHQX1 out_cnt_reg_3_ ( .D(n5836), .CK(clk), .RN(rst_n), .Q(out_cnt[3]) );
  DFFRHQX2 calin_cnt_reg_1_ ( .D(N1363), .CK(clk), .RN(rst_n), .Q(calin_cnt[1]) );
  DFFSX1 out_cnt_6_reg_1_ ( .D(n1719), .CK(clk), .SN(rst_n), .Q(N14321), .QN(
        n727) );
  DFFSX1 out_cnt_6_reg_2_ ( .D(n1721), .CK(clk), .SN(rst_n), .Q(out_cnt_6[2]), 
        .QN(n726) );
  DFFSX1 out_cnt_6_reg_0_ ( .D(n1720), .CK(clk), .SN(rst_n), .Q(out_cnt_6[0]), 
        .QN(n728) );
  DFFRHQX1 c_plus_reg_21_ ( .D(N12587), .CK(clk), .RN(rst_n), .Q(c_plus[21])
         );
  DFFRHQX1 c_plus_reg_17_ ( .D(N12583), .CK(clk), .RN(rst_n), .Q(c_plus[17])
         );
  DFFRHQX1 c_plus_reg_18_ ( .D(N12584), .CK(clk), .RN(rst_n), .Q(c_plus[18])
         );
  DFFRHQX1 c_plus_reg_19_ ( .D(N12585), .CK(clk), .RN(rst_n), .Q(c_plus[19])
         );
  DFFRHQX1 c_plus_reg_24_ ( .D(N12590), .CK(clk), .RN(rst_n), .Q(c_plus[24])
         );
  DFFRHQX1 c_plus_reg_25_ ( .D(N12591), .CK(clk), .RN(rst_n), .Q(c_plus[25])
         );
  DFFRHQX1 c_plus_reg_26_ ( .D(N12592), .CK(clk), .RN(rst_n), .Q(c_plus[26])
         );
  DFFRHQX1 c_plus_reg_29_ ( .D(N12595), .CK(clk), .RN(rst_n), .Q(c_plus[29])
         );
  DFFRHQX1 outset_cnt_reg_3_ ( .D(n1718), .CK(clk), .RN(rst_n), .Q(N945) );
  DFFRHQX1 out_cnt_reg_1_ ( .D(n5838), .CK(clk), .RN(rst_n), .Q(out_cnt[1]) );
  DFFRX1 c_plus_reg_31_ ( .D(N12597), .CK(clk), .RN(rst_n), .QN(n690) );
  DFFRHQX1 c_plus_reg_39_ ( .D(N12605), .CK(clk), .RN(rst_n), .Q(c_plus[39])
         );
  DFFRHQX1 c_plus_reg_33_ ( .D(N12599), .CK(clk), .RN(rst_n), .Q(c_plus[33])
         );
  DFFRHQX1 c_plus_reg_32_ ( .D(N12598), .CK(clk), .RN(rst_n), .Q(c_plus[32])
         );
  DFFRHQX1 c_plus_reg_36_ ( .D(N12602), .CK(clk), .RN(rst_n), .Q(c_plus[36])
         );
  DFFRHQX1 inA11_reg_14_ ( .D(N11408), .CK(clk), .RN(rst_n), .Q(inA11[14]) );
  DFFRHQX1 inA11_reg_15_ ( .D(N11409), .CK(clk), .RN(rst_n), .Q(inA11[15]) );
  DFFRHQX1 w_matrix_reg_0__0__14_ ( .D(n2413), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1022]) );
  DFFRHQX1 w_matrix_reg_0__4__14_ ( .D(n2477), .CK(clk), .RN(rst_n), .Q(
        w_matrix[958]) );
  DFFRHQX1 w_matrix_reg_0__1__14_ ( .D(n2429), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1006]) );
  DFFRHQX1 w_matrix_reg_0__5__14_ ( .D(n2493), .CK(clk), .RN(rst_n), .Q(
        w_matrix[942]) );
  DFFRHQX1 w_matrix_reg_0__2__14_ ( .D(n2445), .CK(clk), .RN(rst_n), .Q(
        w_matrix[990]) );
  DFFRHQX1 w_matrix_reg_0__6__14_ ( .D(n2509), .CK(clk), .RN(rst_n), .Q(
        w_matrix[926]) );
  DFFRHQX1 w_matrix_reg_0__3__14_ ( .D(n2461), .CK(clk), .RN(rst_n), .Q(
        w_matrix[974]) );
  DFFRHQX1 w_matrix_reg_0__7__14_ ( .D(n2525), .CK(clk), .RN(rst_n), .Q(
        w_matrix[910]) );
  DFFRHQX1 w_matrix_reg_0__0__15_ ( .D(n2412), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1023]) );
  DFFRHQX1 w_matrix_reg_0__4__15_ ( .D(n2476), .CK(clk), .RN(rst_n), .Q(
        w_matrix[959]) );
  DFFRHQX1 w_matrix_reg_0__0__13_ ( .D(n2414), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1021]) );
  DFFRHQX1 w_matrix_reg_0__4__13_ ( .D(n2478), .CK(clk), .RN(rst_n), .Q(
        w_matrix[957]) );
  DFFRHQX1 w_matrix_reg_0__0__11_ ( .D(n2416), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1019]) );
  DFFRHQX1 w_matrix_reg_0__4__11_ ( .D(n2480), .CK(clk), .RN(rst_n), .Q(
        w_matrix[955]) );
  DFFRHQX1 w_matrix_reg_0__1__15_ ( .D(n2428), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1007]) );
  DFFRHQX1 w_matrix_reg_0__5__15_ ( .D(n2492), .CK(clk), .RN(rst_n), .Q(
        w_matrix[943]) );
  DFFRHQX1 w_matrix_reg_0__1__13_ ( .D(n2430), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1005]) );
  DFFRHQX1 w_matrix_reg_0__5__13_ ( .D(n2494), .CK(clk), .RN(rst_n), .Q(
        w_matrix[941]) );
  DFFRHQX1 w_matrix_reg_0__1__11_ ( .D(n2432), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1003]) );
  DFFRHQX1 w_matrix_reg_0__5__11_ ( .D(n2496), .CK(clk), .RN(rst_n), .Q(
        w_matrix[939]) );
  DFFRHQX1 w_matrix_reg_0__2__15_ ( .D(n2444), .CK(clk), .RN(rst_n), .Q(
        w_matrix[991]) );
  DFFRHQX1 w_matrix_reg_0__6__15_ ( .D(n2508), .CK(clk), .RN(rst_n), .Q(
        w_matrix[927]) );
  DFFRHQX1 w_matrix_reg_0__2__13_ ( .D(n2446), .CK(clk), .RN(rst_n), .Q(
        w_matrix[989]) );
  DFFRHQX1 w_matrix_reg_0__6__13_ ( .D(n2510), .CK(clk), .RN(rst_n), .Q(
        w_matrix[925]) );
  DFFRHQX1 w_matrix_reg_0__2__11_ ( .D(n2448), .CK(clk), .RN(rst_n), .Q(
        w_matrix[987]) );
  DFFRHQX1 w_matrix_reg_0__6__11_ ( .D(n2512), .CK(clk), .RN(rst_n), .Q(
        w_matrix[923]) );
  DFFRHQX1 w_matrix_reg_0__3__15_ ( .D(n2460), .CK(clk), .RN(rst_n), .Q(
        w_matrix[975]) );
  DFFRHQX1 w_matrix_reg_0__7__15_ ( .D(n2524), .CK(clk), .RN(rst_n), .Q(
        w_matrix[911]) );
  DFFRHQX1 w_matrix_reg_0__3__13_ ( .D(n2462), .CK(clk), .RN(rst_n), .Q(
        w_matrix[973]) );
  DFFRHQX1 w_matrix_reg_0__7__13_ ( .D(n2526), .CK(clk), .RN(rst_n), .Q(
        w_matrix[909]) );
  DFFRHQX1 w_matrix_reg_0__3__11_ ( .D(n2464), .CK(clk), .RN(rst_n), .Q(
        w_matrix[971]) );
  DFFRHQX1 w_matrix_reg_0__7__11_ ( .D(n2528), .CK(clk), .RN(rst_n), .Q(
        w_matrix[907]) );
  DFFRHQX1 inA11_reg_12_ ( .D(N11406), .CK(clk), .RN(rst_n), .Q(inA11[12]) );
  DFFRHQX1 inA11_reg_10_ ( .D(N11404), .CK(clk), .RN(rst_n), .Q(inA11[10]) );
  DFFRHQX1 inA11_reg_8_ ( .D(N11402), .CK(clk), .RN(rst_n), .Q(inA11[8]) );
  DFFRHQX1 inA11_reg_13_ ( .D(N11407), .CK(clk), .RN(rst_n), .Q(inA11[13]) );
  DFFRHQX1 inA11_reg_11_ ( .D(N11405), .CK(clk), .RN(rst_n), .Q(inA11[11]) );
  DFFRHQX1 w_matrix_reg_0__3__9_ ( .D(n2466), .CK(clk), .RN(rst_n), .Q(
        w_matrix[969]) );
  DFFRHQX1 w_matrix_reg_0__7__9_ ( .D(n2530), .CK(clk), .RN(rst_n), .Q(
        w_matrix[905]) );
  DFFRHQX1 w_matrix_reg_0__3__8_ ( .D(n2467), .CK(clk), .RN(rst_n), .Q(
        w_matrix[968]) );
  DFFRHQX1 w_matrix_reg_0__7__8_ ( .D(n2531), .CK(clk), .RN(rst_n), .Q(
        w_matrix[904]) );
  DFFRHQX1 w_matrix_reg_1__4__15_ ( .D(n2604), .CK(clk), .RN(rst_n), .Q(
        w_matrix[831]) );
  DFFRHQX1 w_matrix_reg_2__0__15_ ( .D(n2668), .CK(clk), .RN(rst_n), .Q(
        w_matrix[767]) );
  DFFRHQX1 w_matrix_reg_2__4__15_ ( .D(n2732), .CK(clk), .RN(rst_n), .Q(
        w_matrix[703]) );
  DFFRHQX1 w_matrix_reg_3__0__15_ ( .D(n2796), .CK(clk), .RN(rst_n), .Q(
        w_matrix[639]) );
  DFFRHQX1 w_matrix_reg_3__4__15_ ( .D(n2860), .CK(clk), .RN(rst_n), .Q(
        w_matrix[575]) );
  DFFRHQX1 w_matrix_reg_4__0__15_ ( .D(n2924), .CK(clk), .RN(rst_n), .Q(
        w_matrix[511]) );
  DFFRHQX1 w_matrix_reg_4__4__15_ ( .D(n2988), .CK(clk), .RN(rst_n), .Q(
        w_matrix[447]) );
  DFFRHQX1 w_matrix_reg_5__0__15_ ( .D(n3052), .CK(clk), .RN(rst_n), .Q(
        w_matrix[383]) );
  DFFRHQX1 w_matrix_reg_5__4__15_ ( .D(n3116), .CK(clk), .RN(rst_n), .Q(
        w_matrix[319]) );
  DFFRHQX1 w_matrix_reg_6__0__15_ ( .D(n3180), .CK(clk), .RN(rst_n), .Q(
        w_matrix[255]) );
  DFFRHQX1 w_matrix_reg_6__4__15_ ( .D(n3244), .CK(clk), .RN(rst_n), .Q(
        w_matrix[191]) );
  DFFRHQX1 w_matrix_reg_7__0__15_ ( .D(n3308), .CK(clk), .RN(rst_n), .Q(
        w_matrix[127]) );
  DFFRHQX1 w_matrix_reg_7__4__15_ ( .D(n3372), .CK(clk), .RN(rst_n), .Q(
        w_matrix[63]) );
  DFFRHQX1 w_matrix_reg_0__0__12_ ( .D(n2415), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1020]) );
  DFFRHQX1 w_matrix_reg_0__4__12_ ( .D(n2479), .CK(clk), .RN(rst_n), .Q(
        w_matrix[956]) );
  DFFRHQX1 w_matrix_reg_0__0__10_ ( .D(n2417), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1018]) );
  DFFRHQX1 w_matrix_reg_0__4__10_ ( .D(n2481), .CK(clk), .RN(rst_n), .Q(
        w_matrix[954]) );
  DFFRHQX1 w_matrix_reg_0__0__9_ ( .D(n2418), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1017]) );
  DFFRHQX1 w_matrix_reg_0__4__9_ ( .D(n2482), .CK(clk), .RN(rst_n), .Q(
        w_matrix[953]) );
  DFFRHQX1 w_matrix_reg_0__0__8_ ( .D(n2419), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1016]) );
  DFFRHQX1 w_matrix_reg_0__4__8_ ( .D(n2483), .CK(clk), .RN(rst_n), .Q(
        w_matrix[952]) );
  DFFRHQX1 w_matrix_reg_1__5__15_ ( .D(n2620), .CK(clk), .RN(rst_n), .Q(
        w_matrix[815]) );
  DFFRHQX1 w_matrix_reg_2__1__15_ ( .D(n2684), .CK(clk), .RN(rst_n), .Q(
        w_matrix[751]) );
  DFFRHQX1 w_matrix_reg_2__5__15_ ( .D(n2748), .CK(clk), .RN(rst_n), .Q(
        w_matrix[687]) );
  DFFRHQX1 w_matrix_reg_3__1__15_ ( .D(n2812), .CK(clk), .RN(rst_n), .Q(
        w_matrix[623]) );
  DFFRHQX1 w_matrix_reg_3__5__15_ ( .D(n2876), .CK(clk), .RN(rst_n), .Q(
        w_matrix[559]) );
  DFFRHQX1 w_matrix_reg_4__1__15_ ( .D(n2940), .CK(clk), .RN(rst_n), .Q(
        w_matrix[495]) );
  DFFRHQX1 w_matrix_reg_4__5__15_ ( .D(n3004), .CK(clk), .RN(rst_n), .Q(
        w_matrix[431]) );
  DFFRHQX1 w_matrix_reg_5__1__15_ ( .D(n3068), .CK(clk), .RN(rst_n), .Q(
        w_matrix[367]) );
  DFFRHQX1 w_matrix_reg_5__5__15_ ( .D(n3132), .CK(clk), .RN(rst_n), .Q(
        w_matrix[303]) );
  DFFRHQX1 w_matrix_reg_6__1__15_ ( .D(n3196), .CK(clk), .RN(rst_n), .Q(
        w_matrix[239]) );
  DFFRHQX1 w_matrix_reg_6__5__15_ ( .D(n3260), .CK(clk), .RN(rst_n), .Q(
        w_matrix[175]) );
  DFFRHQX1 w_matrix_reg_7__1__15_ ( .D(n3324), .CK(clk), .RN(rst_n), .Q(
        w_matrix[111]) );
  DFFRHQX1 w_matrix_reg_7__5__15_ ( .D(n3388), .CK(clk), .RN(rst_n), .Q(
        w_matrix[47]) );
  DFFRHQX1 w_matrix_reg_0__1__12_ ( .D(n2431), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1004]) );
  DFFRHQX1 w_matrix_reg_0__5__12_ ( .D(n2495), .CK(clk), .RN(rst_n), .Q(
        w_matrix[940]) );
  DFFRHQX1 w_matrix_reg_0__1__10_ ( .D(n2433), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1002]) );
  DFFRHQX1 w_matrix_reg_0__5__10_ ( .D(n2497), .CK(clk), .RN(rst_n), .Q(
        w_matrix[938]) );
  DFFRHQX1 w_matrix_reg_0__1__9_ ( .D(n2434), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1001]) );
  DFFRHQX1 w_matrix_reg_0__5__9_ ( .D(n2498), .CK(clk), .RN(rst_n), .Q(
        w_matrix[937]) );
  DFFRHQX1 w_matrix_reg_0__1__8_ ( .D(n2435), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1000]) );
  DFFRHQX1 w_matrix_reg_0__5__8_ ( .D(n2499), .CK(clk), .RN(rst_n), .Q(
        w_matrix[936]) );
  DFFRHQX1 w_matrix_reg_1__2__15_ ( .D(n2572), .CK(clk), .RN(rst_n), .Q(
        w_matrix[863]) );
  DFFRHQX1 w_matrix_reg_1__6__15_ ( .D(n2636), .CK(clk), .RN(rst_n), .Q(
        w_matrix[799]) );
  DFFRHQX1 w_matrix_reg_2__2__15_ ( .D(n2700), .CK(clk), .RN(rst_n), .Q(
        w_matrix[735]) );
  DFFRHQX1 w_matrix_reg_2__6__15_ ( .D(n2764), .CK(clk), .RN(rst_n), .Q(
        w_matrix[671]) );
  DFFRHQX1 w_matrix_reg_3__2__15_ ( .D(n2828), .CK(clk), .RN(rst_n), .Q(
        w_matrix[607]) );
  DFFRHQX1 w_matrix_reg_3__6__15_ ( .D(n2892), .CK(clk), .RN(rst_n), .Q(
        w_matrix[543]) );
  DFFRHQX1 w_matrix_reg_4__2__15_ ( .D(n2956), .CK(clk), .RN(rst_n), .Q(
        w_matrix[479]) );
  DFFRHQX1 w_matrix_reg_4__6__15_ ( .D(n3020), .CK(clk), .RN(rst_n), .Q(
        w_matrix[415]) );
  DFFRHQX1 w_matrix_reg_5__2__15_ ( .D(n3084), .CK(clk), .RN(rst_n), .Q(
        w_matrix[351]) );
  DFFRHQX1 w_matrix_reg_5__6__15_ ( .D(n3148), .CK(clk), .RN(rst_n), .Q(
        w_matrix[287]) );
  DFFRHQX1 w_matrix_reg_6__2__15_ ( .D(n3212), .CK(clk), .RN(rst_n), .Q(
        w_matrix[223]) );
  DFFRHQX1 w_matrix_reg_6__6__15_ ( .D(n3276), .CK(clk), .RN(rst_n), .Q(
        w_matrix[159]) );
  DFFRHQX1 w_matrix_reg_7__2__15_ ( .D(n3340), .CK(clk), .RN(rst_n), .Q(
        w_matrix[95]) );
  DFFRHQX1 w_matrix_reg_7__6__15_ ( .D(n3404), .CK(clk), .RN(rst_n), .Q(
        w_matrix[31]) );
  DFFRHQX1 w_matrix_reg_0__2__12_ ( .D(n2447), .CK(clk), .RN(rst_n), .Q(
        w_matrix[988]) );
  DFFRHQX1 w_matrix_reg_0__6__12_ ( .D(n2511), .CK(clk), .RN(rst_n), .Q(
        w_matrix[924]) );
  DFFRHQX1 w_matrix_reg_0__2__10_ ( .D(n2449), .CK(clk), .RN(rst_n), .Q(
        w_matrix[986]) );
  DFFRHQX1 w_matrix_reg_0__6__10_ ( .D(n2513), .CK(clk), .RN(rst_n), .Q(
        w_matrix[922]) );
  DFFRHQX1 w_matrix_reg_0__2__9_ ( .D(n2450), .CK(clk), .RN(rst_n), .Q(
        w_matrix[985]) );
  DFFRHQX1 w_matrix_reg_0__6__9_ ( .D(n2514), .CK(clk), .RN(rst_n), .Q(
        w_matrix[921]) );
  DFFRHQX1 w_matrix_reg_0__2__8_ ( .D(n2451), .CK(clk), .RN(rst_n), .Q(
        w_matrix[984]) );
  DFFRHQX1 w_matrix_reg_0__6__8_ ( .D(n2515), .CK(clk), .RN(rst_n), .Q(
        w_matrix[920]) );
  DFFRHQX1 w_matrix_reg_1__3__15_ ( .D(n2588), .CK(clk), .RN(rst_n), .Q(
        w_matrix[847]) );
  DFFRHQX1 w_matrix_reg_1__7__15_ ( .D(n2652), .CK(clk), .RN(rst_n), .Q(
        w_matrix[783]) );
  DFFRHQX1 w_matrix_reg_2__3__15_ ( .D(n2716), .CK(clk), .RN(rst_n), .Q(
        w_matrix[719]) );
  DFFRHQX1 w_matrix_reg_2__7__15_ ( .D(n2780), .CK(clk), .RN(rst_n), .Q(
        w_matrix[655]) );
  DFFRHQX1 w_matrix_reg_3__3__15_ ( .D(n2844), .CK(clk), .RN(rst_n), .Q(
        w_matrix[591]) );
  DFFRHQX1 w_matrix_reg_3__7__15_ ( .D(n2908), .CK(clk), .RN(rst_n), .Q(
        w_matrix[527]) );
  DFFRHQX1 w_matrix_reg_4__3__15_ ( .D(n2972), .CK(clk), .RN(rst_n), .Q(
        w_matrix[463]) );
  DFFRHQX1 w_matrix_reg_4__7__15_ ( .D(n3036), .CK(clk), .RN(rst_n), .Q(
        w_matrix[399]) );
  DFFRHQX1 w_matrix_reg_5__3__15_ ( .D(n3100), .CK(clk), .RN(rst_n), .Q(
        w_matrix[335]) );
  DFFRHQX1 w_matrix_reg_5__7__15_ ( .D(n3164), .CK(clk), .RN(rst_n), .Q(
        w_matrix[271]) );
  DFFRHQX1 w_matrix_reg_6__3__15_ ( .D(n3228), .CK(clk), .RN(rst_n), .Q(
        w_matrix[207]) );
  DFFRHQX1 w_matrix_reg_6__7__15_ ( .D(n3292), .CK(clk), .RN(rst_n), .Q(
        w_matrix[143]) );
  DFFRHQX1 w_matrix_reg_7__3__15_ ( .D(n3356), .CK(clk), .RN(rst_n), .Q(
        w_matrix[79]) );
  DFFRHQX1 w_matrix_reg_7__7__15_ ( .D(n3420), .CK(clk), .RN(rst_n), .Q(
        w_matrix[15]) );
  DFFRHQX1 w_matrix_reg_0__3__12_ ( .D(n2463), .CK(clk), .RN(rst_n), .Q(
        w_matrix[972]) );
  DFFRHQX1 w_matrix_reg_0__7__12_ ( .D(n2527), .CK(clk), .RN(rst_n), .Q(
        w_matrix[908]) );
  DFFRHQX1 w_matrix_reg_0__3__10_ ( .D(n2465), .CK(clk), .RN(rst_n), .Q(
        w_matrix[970]) );
  DFFRHQX1 w_matrix_reg_0__7__10_ ( .D(n2529), .CK(clk), .RN(rst_n), .Q(
        w_matrix[906]) );
  DFFRX1 w_matrix_reg_1__1__14_ ( .D(n2557), .CK(clk), .RN(rst_n), .Q(
        w_matrix[878]), .QN(n659) );
  DFFRX1 w_matrix_reg_1__1__15_ ( .D(n2556), .CK(clk), .RN(rst_n), .Q(
        w_matrix[879]), .QN(n658) );
  DFFRX1 w_matrix_reg_1__1__13_ ( .D(n2558), .CK(clk), .RN(rst_n), .Q(
        w_matrix[877]), .QN(n660) );
  DFFRHQX1 inA51_reg_14_ ( .D(N11787), .CK(clk), .RN(rst_n), .Q(inA51[14]) );
  DFFRHQX1 inA51_reg_12_ ( .D(N11785), .CK(clk), .RN(rst_n), .Q(inA51[12]) );
  DFFRHQX1 inA61_reg_14_ ( .D(N11884), .CK(clk), .RN(rst_n), .Q(inA61[14]) );
  DFFRHQX1 inA61_reg_12_ ( .D(N11882), .CK(clk), .RN(rst_n), .Q(inA61[12]) );
  DFFRHQX1 inA31_reg_14_ ( .D(N11598), .CK(clk), .RN(rst_n), .Q(inA31[14]) );
  DFFRHQX1 inA71_reg_14_ ( .D(N11978), .CK(clk), .RN(rst_n), .Q(inA71[14]) );
  DFFRHQX1 inA31_reg_12_ ( .D(N11596), .CK(clk), .RN(rst_n), .Q(inA31[12]) );
  DFFRHQX1 inA71_reg_12_ ( .D(N11976), .CK(clk), .RN(rst_n), .Q(inA71[12]) );
  DFFRHQX1 inA11_reg_6_ ( .D(N11400), .CK(clk), .RN(rst_n), .Q(inA11[6]) );
  DFFRHQX1 inA11_reg_4_ ( .D(N11398), .CK(clk), .RN(rst_n), .Q(inA11[4]) );
  DFFRHQX1 inA11_reg_2_ ( .D(N11396), .CK(clk), .RN(rst_n), .Q(inA11[2]) );
  DFFRHQX1 inA21_reg_14_ ( .D(N11504), .CK(clk), .RN(rst_n), .Q(inA21[14]) );
  DFFRHQX1 inA41_reg_14_ ( .D(N11695), .CK(clk), .RN(rst_n), .Q(inA41[14]) );
  DFFRHQX1 inA81_reg_14_ ( .D(N12074), .CK(clk), .RN(rst_n), .Q(inA81[14]) );
  DFFRHQX1 inA21_reg_12_ ( .D(N11502), .CK(clk), .RN(rst_n), .Q(inA21[12]) );
  DFFRHQX1 inA41_reg_12_ ( .D(N11693), .CK(clk), .RN(rst_n), .Q(inA41[12]) );
  DFFRHQX1 inA81_reg_12_ ( .D(N12072), .CK(clk), .RN(rst_n), .Q(inA81[12]) );
  DFFRHQX1 inA51_reg_15_ ( .D(N11788), .CK(clk), .RN(rst_n), .Q(inA51[15]) );
  DFFRHQX1 inA61_reg_15_ ( .D(N11885), .CK(clk), .RN(rst_n), .Q(inA61[15]) );
  DFFRHQX1 inA31_reg_15_ ( .D(N11599), .CK(clk), .RN(rst_n), .Q(inA31[15]) );
  DFFRHQX1 inA71_reg_15_ ( .D(N11979), .CK(clk), .RN(rst_n), .Q(inA71[15]) );
  DFFRHQX1 inA11_reg_9_ ( .D(N11403), .CK(clk), .RN(rst_n), .Q(inA11[9]) );
  DFFRHQX1 inA11_reg_7_ ( .D(N11401), .CK(clk), .RN(rst_n), .Q(inA11[7]) );
  DFFRHQX1 inA11_reg_5_ ( .D(N11399), .CK(clk), .RN(rst_n), .Q(inA11[5]) );
  DFFRHQX1 inA21_reg_15_ ( .D(N11505), .CK(clk), .RN(rst_n), .Q(inA21[15]) );
  DFFRHQX1 inA41_reg_15_ ( .D(N11696), .CK(clk), .RN(rst_n), .Q(inA41[15]) );
  DFFRHQX1 inA81_reg_15_ ( .D(N12075), .CK(clk), .RN(rst_n), .Q(inA81[15]) );
  DFFRHQX1 w_matrix_reg_0__0__0_ ( .D(n2427), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1008]) );
  DFFRHQX1 w_matrix_reg_0__4__0_ ( .D(n2491), .CK(clk), .RN(rst_n), .Q(
        w_matrix[944]) );
  DFFRHQX1 w_matrix_reg_0__1__0_ ( .D(n2443), .CK(clk), .RN(rst_n), .Q(
        w_matrix[992]) );
  DFFRHQX1 w_matrix_reg_0__5__0_ ( .D(n2507), .CK(clk), .RN(rst_n), .Q(
        w_matrix[928]) );
  DFFRHQX1 w_matrix_reg_0__2__0_ ( .D(n2459), .CK(clk), .RN(rst_n), .Q(
        w_matrix[976]) );
  DFFRHQX1 w_matrix_reg_0__6__0_ ( .D(n2523), .CK(clk), .RN(rst_n), .Q(
        w_matrix[912]) );
  DFFRHQX1 w_matrix_reg_0__3__0_ ( .D(n2475), .CK(clk), .RN(rst_n), .Q(
        w_matrix[960]) );
  DFFRHQX1 w_matrix_reg_0__7__0_ ( .D(n2539), .CK(clk), .RN(rst_n), .Q(
        w_matrix[896]) );
  DFFRHQX1 w_matrix_reg_1__4__14_ ( .D(n2605), .CK(clk), .RN(rst_n), .Q(
        w_matrix[830]) );
  DFFRHQX1 w_matrix_reg_2__0__14_ ( .D(n2669), .CK(clk), .RN(rst_n), .Q(
        w_matrix[766]) );
  DFFRHQX1 w_matrix_reg_2__4__14_ ( .D(n2733), .CK(clk), .RN(rst_n), .Q(
        w_matrix[702]) );
  DFFRHQX1 w_matrix_reg_3__0__14_ ( .D(n2797), .CK(clk), .RN(rst_n), .Q(
        w_matrix[638]) );
  DFFRHQX1 w_matrix_reg_3__4__14_ ( .D(n2861), .CK(clk), .RN(rst_n), .Q(
        w_matrix[574]) );
  DFFRHQX1 w_matrix_reg_4__0__14_ ( .D(n2925), .CK(clk), .RN(rst_n), .Q(
        w_matrix[510]) );
  DFFRHQX1 w_matrix_reg_4__4__14_ ( .D(n2989), .CK(clk), .RN(rst_n), .Q(
        w_matrix[446]) );
  DFFRHQX1 w_matrix_reg_5__0__14_ ( .D(n3053), .CK(clk), .RN(rst_n), .Q(
        w_matrix[382]) );
  DFFRHQX1 w_matrix_reg_5__4__14_ ( .D(n3117), .CK(clk), .RN(rst_n), .Q(
        w_matrix[318]) );
  DFFRHQX1 w_matrix_reg_6__0__14_ ( .D(n3181), .CK(clk), .RN(rst_n), .Q(
        w_matrix[254]) );
  DFFRHQX1 w_matrix_reg_6__4__14_ ( .D(n3245), .CK(clk), .RN(rst_n), .Q(
        w_matrix[190]) );
  DFFRHQX1 w_matrix_reg_7__0__14_ ( .D(n3309), .CK(clk), .RN(rst_n), .Q(
        w_matrix[126]) );
  DFFRHQX1 w_matrix_reg_7__4__14_ ( .D(n3373), .CK(clk), .RN(rst_n), .Q(
        w_matrix[62]) );
  DFFRHQX1 w_matrix_reg_1__5__14_ ( .D(n2621), .CK(clk), .RN(rst_n), .Q(
        w_matrix[814]) );
  DFFRHQX1 w_matrix_reg_2__1__14_ ( .D(n2685), .CK(clk), .RN(rst_n), .Q(
        w_matrix[750]) );
  DFFRHQX1 w_matrix_reg_2__5__14_ ( .D(n2749), .CK(clk), .RN(rst_n), .Q(
        w_matrix[686]) );
  DFFRHQX1 w_matrix_reg_3__1__14_ ( .D(n2813), .CK(clk), .RN(rst_n), .Q(
        w_matrix[622]) );
  DFFRHQX1 w_matrix_reg_3__5__14_ ( .D(n2877), .CK(clk), .RN(rst_n), .Q(
        w_matrix[558]) );
  DFFRHQX1 w_matrix_reg_4__1__14_ ( .D(n2941), .CK(clk), .RN(rst_n), .Q(
        w_matrix[494]) );
  DFFRHQX1 w_matrix_reg_4__5__14_ ( .D(n3005), .CK(clk), .RN(rst_n), .Q(
        w_matrix[430]) );
  DFFRHQX1 w_matrix_reg_5__1__14_ ( .D(n3069), .CK(clk), .RN(rst_n), .Q(
        w_matrix[366]) );
  DFFRHQX1 w_matrix_reg_5__5__14_ ( .D(n3133), .CK(clk), .RN(rst_n), .Q(
        w_matrix[302]) );
  DFFRHQX1 w_matrix_reg_6__1__14_ ( .D(n3197), .CK(clk), .RN(rst_n), .Q(
        w_matrix[238]) );
  DFFRHQX1 w_matrix_reg_6__5__14_ ( .D(n3261), .CK(clk), .RN(rst_n), .Q(
        w_matrix[174]) );
  DFFRHQX1 w_matrix_reg_7__1__14_ ( .D(n3325), .CK(clk), .RN(rst_n), .Q(
        w_matrix[110]) );
  DFFRHQX1 w_matrix_reg_7__5__14_ ( .D(n3389), .CK(clk), .RN(rst_n), .Q(
        w_matrix[46]) );
  DFFRHQX1 w_matrix_reg_1__2__14_ ( .D(n2573), .CK(clk), .RN(rst_n), .Q(
        w_matrix[862]) );
  DFFRHQX1 w_matrix_reg_1__6__14_ ( .D(n2637), .CK(clk), .RN(rst_n), .Q(
        w_matrix[798]) );
  DFFRHQX1 w_matrix_reg_2__2__14_ ( .D(n2701), .CK(clk), .RN(rst_n), .Q(
        w_matrix[734]) );
  DFFRHQX1 w_matrix_reg_2__6__14_ ( .D(n2765), .CK(clk), .RN(rst_n), .Q(
        w_matrix[670]) );
  DFFRHQX1 w_matrix_reg_3__2__14_ ( .D(n2829), .CK(clk), .RN(rst_n), .Q(
        w_matrix[606]) );
  DFFRHQX1 w_matrix_reg_3__6__14_ ( .D(n2893), .CK(clk), .RN(rst_n), .Q(
        w_matrix[542]) );
  DFFRHQX1 w_matrix_reg_4__2__14_ ( .D(n2957), .CK(clk), .RN(rst_n), .Q(
        w_matrix[478]) );
  DFFRHQX1 w_matrix_reg_4__6__14_ ( .D(n3021), .CK(clk), .RN(rst_n), .Q(
        w_matrix[414]) );
  DFFRHQX1 w_matrix_reg_5__2__14_ ( .D(n3085), .CK(clk), .RN(rst_n), .Q(
        w_matrix[350]) );
  DFFRHQX1 w_matrix_reg_5__6__14_ ( .D(n3149), .CK(clk), .RN(rst_n), .Q(
        w_matrix[286]) );
  DFFRHQX1 w_matrix_reg_6__2__14_ ( .D(n3213), .CK(clk), .RN(rst_n), .Q(
        w_matrix[222]) );
  DFFRHQX1 w_matrix_reg_6__6__14_ ( .D(n3277), .CK(clk), .RN(rst_n), .Q(
        w_matrix[158]) );
  DFFRHQX1 w_matrix_reg_7__2__14_ ( .D(n3341), .CK(clk), .RN(rst_n), .Q(
        w_matrix[94]) );
  DFFRHQX1 w_matrix_reg_7__6__14_ ( .D(n3405), .CK(clk), .RN(rst_n), .Q(
        w_matrix[30]) );
  DFFRHQX1 w_matrix_reg_1__3__14_ ( .D(n2589), .CK(clk), .RN(rst_n), .Q(
        w_matrix[846]) );
  DFFRHQX1 w_matrix_reg_1__7__14_ ( .D(n2653), .CK(clk), .RN(rst_n), .Q(
        w_matrix[782]) );
  DFFRHQX1 w_matrix_reg_2__3__14_ ( .D(n2717), .CK(clk), .RN(rst_n), .Q(
        w_matrix[718]) );
  DFFRHQX1 w_matrix_reg_2__7__14_ ( .D(n2781), .CK(clk), .RN(rst_n), .Q(
        w_matrix[654]) );
  DFFRHQX1 w_matrix_reg_3__3__14_ ( .D(n2845), .CK(clk), .RN(rst_n), .Q(
        w_matrix[590]) );
  DFFRHQX1 w_matrix_reg_3__7__14_ ( .D(n2909), .CK(clk), .RN(rst_n), .Q(
        w_matrix[526]) );
  DFFRHQX1 w_matrix_reg_4__3__14_ ( .D(n2973), .CK(clk), .RN(rst_n), .Q(
        w_matrix[462]) );
  DFFRHQX1 w_matrix_reg_4__7__14_ ( .D(n3037), .CK(clk), .RN(rst_n), .Q(
        w_matrix[398]) );
  DFFRHQX1 w_matrix_reg_5__3__14_ ( .D(n3101), .CK(clk), .RN(rst_n), .Q(
        w_matrix[334]) );
  DFFRHQX1 w_matrix_reg_5__7__14_ ( .D(n3165), .CK(clk), .RN(rst_n), .Q(
        w_matrix[270]) );
  DFFRHQX1 w_matrix_reg_6__3__14_ ( .D(n3229), .CK(clk), .RN(rst_n), .Q(
        w_matrix[206]) );
  DFFRHQX1 w_matrix_reg_6__7__14_ ( .D(n3293), .CK(clk), .RN(rst_n), .Q(
        w_matrix[142]) );
  DFFRHQX1 w_matrix_reg_7__3__14_ ( .D(n3357), .CK(clk), .RN(rst_n), .Q(
        w_matrix[78]) );
  DFFRHQX1 w_matrix_reg_7__7__14_ ( .D(n3421), .CK(clk), .RN(rst_n), .Q(
        w_matrix[14]) );
  DFFRHQX1 w_matrix_reg_0__3__7_ ( .D(n2468), .CK(clk), .RN(rst_n), .Q(
        w_matrix[967]) );
  DFFRHQX1 w_matrix_reg_0__7__7_ ( .D(n2532), .CK(clk), .RN(rst_n), .Q(
        w_matrix[903]) );
  DFFRHQX1 w_matrix_reg_0__3__6_ ( .D(n2469), .CK(clk), .RN(rst_n), .Q(
        w_matrix[966]) );
  DFFRHQX1 w_matrix_reg_0__7__6_ ( .D(n2533), .CK(clk), .RN(rst_n), .Q(
        w_matrix[902]) );
  DFFRHQX1 w_matrix_reg_1__4__13_ ( .D(n2606), .CK(clk), .RN(rst_n), .Q(
        w_matrix[829]) );
  DFFRHQX1 w_matrix_reg_2__0__13_ ( .D(n2670), .CK(clk), .RN(rst_n), .Q(
        w_matrix[765]) );
  DFFRHQX1 w_matrix_reg_2__4__13_ ( .D(n2734), .CK(clk), .RN(rst_n), .Q(
        w_matrix[701]) );
  DFFRHQX1 w_matrix_reg_3__0__13_ ( .D(n2798), .CK(clk), .RN(rst_n), .Q(
        w_matrix[637]) );
  DFFRHQX1 w_matrix_reg_3__4__13_ ( .D(n2862), .CK(clk), .RN(rst_n), .Q(
        w_matrix[573]) );
  DFFRHQX1 w_matrix_reg_4__0__13_ ( .D(n2926), .CK(clk), .RN(rst_n), .Q(
        w_matrix[509]) );
  DFFRHQX1 w_matrix_reg_4__4__13_ ( .D(n2990), .CK(clk), .RN(rst_n), .Q(
        w_matrix[445]) );
  DFFRHQX1 w_matrix_reg_5__0__13_ ( .D(n3054), .CK(clk), .RN(rst_n), .Q(
        w_matrix[381]) );
  DFFRHQX1 w_matrix_reg_5__4__13_ ( .D(n3118), .CK(clk), .RN(rst_n), .Q(
        w_matrix[317]) );
  DFFRHQX1 w_matrix_reg_6__0__13_ ( .D(n3182), .CK(clk), .RN(rst_n), .Q(
        w_matrix[253]) );
  DFFRHQX1 w_matrix_reg_6__4__13_ ( .D(n3246), .CK(clk), .RN(rst_n), .Q(
        w_matrix[189]) );
  DFFRHQX1 w_matrix_reg_7__0__13_ ( .D(n3310), .CK(clk), .RN(rst_n), .Q(
        w_matrix[125]) );
  DFFRHQX1 w_matrix_reg_7__4__13_ ( .D(n3374), .CK(clk), .RN(rst_n), .Q(
        w_matrix[61]) );
  DFFRHQX1 w_matrix_reg_1__4__12_ ( .D(n2607), .CK(clk), .RN(rst_n), .Q(
        w_matrix[828]) );
  DFFRHQX1 w_matrix_reg_2__0__12_ ( .D(n2671), .CK(clk), .RN(rst_n), .Q(
        w_matrix[764]) );
  DFFRHQX1 w_matrix_reg_2__4__12_ ( .D(n2735), .CK(clk), .RN(rst_n), .Q(
        w_matrix[700]) );
  DFFRHQX1 w_matrix_reg_3__0__12_ ( .D(n2799), .CK(clk), .RN(rst_n), .Q(
        w_matrix[636]) );
  DFFRHQX1 w_matrix_reg_3__4__12_ ( .D(n2863), .CK(clk), .RN(rst_n), .Q(
        w_matrix[572]) );
  DFFRHQX1 w_matrix_reg_4__0__12_ ( .D(n2927), .CK(clk), .RN(rst_n), .Q(
        w_matrix[508]) );
  DFFRHQX1 w_matrix_reg_4__4__12_ ( .D(n2991), .CK(clk), .RN(rst_n), .Q(
        w_matrix[444]) );
  DFFRHQX1 w_matrix_reg_5__0__12_ ( .D(n3055), .CK(clk), .RN(rst_n), .Q(
        w_matrix[380]) );
  DFFRHQX1 w_matrix_reg_5__4__12_ ( .D(n3119), .CK(clk), .RN(rst_n), .Q(
        w_matrix[316]) );
  DFFRHQX1 w_matrix_reg_6__0__12_ ( .D(n3183), .CK(clk), .RN(rst_n), .Q(
        w_matrix[252]) );
  DFFRHQX1 w_matrix_reg_6__4__12_ ( .D(n3247), .CK(clk), .RN(rst_n), .Q(
        w_matrix[188]) );
  DFFRHQX1 w_matrix_reg_7__0__12_ ( .D(n3311), .CK(clk), .RN(rst_n), .Q(
        w_matrix[124]) );
  DFFRHQX1 w_matrix_reg_7__4__12_ ( .D(n3375), .CK(clk), .RN(rst_n), .Q(
        w_matrix[60]) );
  DFFRHQX1 w_matrix_reg_0__3__5_ ( .D(n2470), .CK(clk), .RN(rst_n), .Q(
        w_matrix[965]) );
  DFFRHQX1 w_matrix_reg_0__7__5_ ( .D(n2534), .CK(clk), .RN(rst_n), .Q(
        w_matrix[901]) );
  DFFRHQX1 w_matrix_reg_1__4__11_ ( .D(n2608), .CK(clk), .RN(rst_n), .Q(
        w_matrix[827]) );
  DFFRHQX1 w_matrix_reg_2__0__11_ ( .D(n2672), .CK(clk), .RN(rst_n), .Q(
        w_matrix[763]) );
  DFFRHQX1 w_matrix_reg_2__4__11_ ( .D(n2736), .CK(clk), .RN(rst_n), .Q(
        w_matrix[699]) );
  DFFRHQX1 w_matrix_reg_3__0__11_ ( .D(n2800), .CK(clk), .RN(rst_n), .Q(
        w_matrix[635]) );
  DFFRHQX1 w_matrix_reg_3__4__11_ ( .D(n2864), .CK(clk), .RN(rst_n), .Q(
        w_matrix[571]) );
  DFFRHQX1 w_matrix_reg_4__0__11_ ( .D(n2928), .CK(clk), .RN(rst_n), .Q(
        w_matrix[507]) );
  DFFRHQX1 w_matrix_reg_4__4__11_ ( .D(n2992), .CK(clk), .RN(rst_n), .Q(
        w_matrix[443]) );
  DFFRHQX1 w_matrix_reg_5__0__11_ ( .D(n3056), .CK(clk), .RN(rst_n), .Q(
        w_matrix[379]) );
  DFFRHQX1 w_matrix_reg_5__4__11_ ( .D(n3120), .CK(clk), .RN(rst_n), .Q(
        w_matrix[315]) );
  DFFRHQX1 w_matrix_reg_6__0__11_ ( .D(n3184), .CK(clk), .RN(rst_n), .Q(
        w_matrix[251]) );
  DFFRHQX1 w_matrix_reg_6__4__11_ ( .D(n3248), .CK(clk), .RN(rst_n), .Q(
        w_matrix[187]) );
  DFFRHQX1 w_matrix_reg_7__0__11_ ( .D(n3312), .CK(clk), .RN(rst_n), .Q(
        w_matrix[123]) );
  DFFRHQX1 w_matrix_reg_7__4__11_ ( .D(n3376), .CK(clk), .RN(rst_n), .Q(
        w_matrix[59]) );
  DFFRHQX1 w_matrix_reg_0__0__7_ ( .D(n2420), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1015]) );
  DFFRHQX1 w_matrix_reg_0__4__7_ ( .D(n2484), .CK(clk), .RN(rst_n), .Q(
        w_matrix[951]) );
  DFFRHQX1 w_matrix_reg_0__0__6_ ( .D(n2421), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1014]) );
  DFFRHQX1 w_matrix_reg_0__4__6_ ( .D(n2485), .CK(clk), .RN(rst_n), .Q(
        w_matrix[950]) );
  DFFRHQX1 w_matrix_reg_0__0__5_ ( .D(n2422), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1013]) );
  DFFRHQX1 w_matrix_reg_0__4__5_ ( .D(n2486), .CK(clk), .RN(rst_n), .Q(
        w_matrix[949]) );
  DFFRHQX1 w_matrix_reg_0__0__4_ ( .D(n2423), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1012]) );
  DFFRHQX1 w_matrix_reg_0__4__4_ ( .D(n2487), .CK(clk), .RN(rst_n), .Q(
        w_matrix[948]) );
  DFFRHQX1 w_matrix_reg_0__0__3_ ( .D(n2424), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1011]) );
  DFFRHQX1 w_matrix_reg_0__4__3_ ( .D(n2488), .CK(clk), .RN(rst_n), .Q(
        w_matrix[947]) );
  DFFRHQX1 w_matrix_reg_0__0__2_ ( .D(n2425), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1010]) );
  DFFRHQX1 w_matrix_reg_0__4__2_ ( .D(n2489), .CK(clk), .RN(rst_n), .Q(
        w_matrix[946]) );
  DFFRHQX1 w_matrix_reg_0__3__4_ ( .D(n2471), .CK(clk), .RN(rst_n), .Q(
        w_matrix[964]) );
  DFFRHQX1 w_matrix_reg_0__7__4_ ( .D(n2535), .CK(clk), .RN(rst_n), .Q(
        w_matrix[900]) );
  DFFRHQX1 w_matrix_reg_0__0__1_ ( .D(n2426), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1009]) );
  DFFRHQX1 w_matrix_reg_0__4__1_ ( .D(n2490), .CK(clk), .RN(rst_n), .Q(
        w_matrix[945]) );
  DFFRHQX1 w_matrix_reg_1__5__13_ ( .D(n2622), .CK(clk), .RN(rst_n), .Q(
        w_matrix[813]) );
  DFFRHQX1 w_matrix_reg_2__1__13_ ( .D(n2686), .CK(clk), .RN(rst_n), .Q(
        w_matrix[749]) );
  DFFRHQX1 w_matrix_reg_2__5__13_ ( .D(n2750), .CK(clk), .RN(rst_n), .Q(
        w_matrix[685]) );
  DFFRHQX1 w_matrix_reg_3__1__13_ ( .D(n2814), .CK(clk), .RN(rst_n), .Q(
        w_matrix[621]) );
  DFFRHQX1 w_matrix_reg_3__5__13_ ( .D(n2878), .CK(clk), .RN(rst_n), .Q(
        w_matrix[557]) );
  DFFRHQX1 w_matrix_reg_4__1__13_ ( .D(n2942), .CK(clk), .RN(rst_n), .Q(
        w_matrix[493]) );
  DFFRHQX1 w_matrix_reg_4__5__13_ ( .D(n3006), .CK(clk), .RN(rst_n), .Q(
        w_matrix[429]) );
  DFFRHQX1 w_matrix_reg_5__1__13_ ( .D(n3070), .CK(clk), .RN(rst_n), .Q(
        w_matrix[365]) );
  DFFRHQX1 w_matrix_reg_5__5__13_ ( .D(n3134), .CK(clk), .RN(rst_n), .Q(
        w_matrix[301]) );
  DFFRHQX1 w_matrix_reg_6__1__13_ ( .D(n3198), .CK(clk), .RN(rst_n), .Q(
        w_matrix[237]) );
  DFFRHQX1 w_matrix_reg_6__5__13_ ( .D(n3262), .CK(clk), .RN(rst_n), .Q(
        w_matrix[173]) );
  DFFRHQX1 w_matrix_reg_7__1__13_ ( .D(n3326), .CK(clk), .RN(rst_n), .Q(
        w_matrix[109]) );
  DFFRHQX1 w_matrix_reg_7__5__13_ ( .D(n3390), .CK(clk), .RN(rst_n), .Q(
        w_matrix[45]) );
  DFFRHQX1 w_matrix_reg_1__5__12_ ( .D(n2623), .CK(clk), .RN(rst_n), .Q(
        w_matrix[812]) );
  DFFRHQX1 w_matrix_reg_2__1__12_ ( .D(n2687), .CK(clk), .RN(rst_n), .Q(
        w_matrix[748]) );
  DFFRHQX1 w_matrix_reg_2__5__12_ ( .D(n2751), .CK(clk), .RN(rst_n), .Q(
        w_matrix[684]) );
  DFFRHQX1 w_matrix_reg_3__1__12_ ( .D(n2815), .CK(clk), .RN(rst_n), .Q(
        w_matrix[620]) );
  DFFRHQX1 w_matrix_reg_3__5__12_ ( .D(n2879), .CK(clk), .RN(rst_n), .Q(
        w_matrix[556]) );
  DFFRHQX1 w_matrix_reg_4__1__12_ ( .D(n2943), .CK(clk), .RN(rst_n), .Q(
        w_matrix[492]) );
  DFFRHQX1 w_matrix_reg_4__5__12_ ( .D(n3007), .CK(clk), .RN(rst_n), .Q(
        w_matrix[428]) );
  DFFRHQX1 w_matrix_reg_5__1__12_ ( .D(n3071), .CK(clk), .RN(rst_n), .Q(
        w_matrix[364]) );
  DFFRHQX1 w_matrix_reg_5__5__12_ ( .D(n3135), .CK(clk), .RN(rst_n), .Q(
        w_matrix[300]) );
  DFFRHQX1 w_matrix_reg_6__1__12_ ( .D(n3199), .CK(clk), .RN(rst_n), .Q(
        w_matrix[236]) );
  DFFRHQX1 w_matrix_reg_6__5__12_ ( .D(n3263), .CK(clk), .RN(rst_n), .Q(
        w_matrix[172]) );
  DFFRHQX1 w_matrix_reg_7__1__12_ ( .D(n3327), .CK(clk), .RN(rst_n), .Q(
        w_matrix[108]) );
  DFFRHQX1 w_matrix_reg_7__5__12_ ( .D(n3391), .CK(clk), .RN(rst_n), .Q(
        w_matrix[44]) );
  DFFRHQX1 w_matrix_reg_1__5__11_ ( .D(n2624), .CK(clk), .RN(rst_n), .Q(
        w_matrix[811]) );
  DFFRHQX1 w_matrix_reg_2__1__11_ ( .D(n2688), .CK(clk), .RN(rst_n), .Q(
        w_matrix[747]) );
  DFFRHQX1 w_matrix_reg_2__5__11_ ( .D(n2752), .CK(clk), .RN(rst_n), .Q(
        w_matrix[683]) );
  DFFRHQX1 w_matrix_reg_3__1__11_ ( .D(n2816), .CK(clk), .RN(rst_n), .Q(
        w_matrix[619]) );
  DFFRHQX1 w_matrix_reg_3__5__11_ ( .D(n2880), .CK(clk), .RN(rst_n), .Q(
        w_matrix[555]) );
  DFFRHQX1 w_matrix_reg_4__1__11_ ( .D(n2944), .CK(clk), .RN(rst_n), .Q(
        w_matrix[491]) );
  DFFRHQX1 w_matrix_reg_4__5__11_ ( .D(n3008), .CK(clk), .RN(rst_n), .Q(
        w_matrix[427]) );
  DFFRHQX1 w_matrix_reg_5__1__11_ ( .D(n3072), .CK(clk), .RN(rst_n), .Q(
        w_matrix[363]) );
  DFFRHQX1 w_matrix_reg_5__5__11_ ( .D(n3136), .CK(clk), .RN(rst_n), .Q(
        w_matrix[299]) );
  DFFRHQX1 w_matrix_reg_6__1__11_ ( .D(n3200), .CK(clk), .RN(rst_n), .Q(
        w_matrix[235]) );
  DFFRHQX1 w_matrix_reg_6__5__11_ ( .D(n3264), .CK(clk), .RN(rst_n), .Q(
        w_matrix[171]) );
  DFFRHQX1 w_matrix_reg_7__1__11_ ( .D(n3328), .CK(clk), .RN(rst_n), .Q(
        w_matrix[107]) );
  DFFRHQX1 w_matrix_reg_7__5__11_ ( .D(n3392), .CK(clk), .RN(rst_n), .Q(
        w_matrix[43]) );
  DFFRHQX1 w_matrix_reg_0__3__3_ ( .D(n2472), .CK(clk), .RN(rst_n), .Q(
        w_matrix[963]) );
  DFFRHQX1 w_matrix_reg_0__7__3_ ( .D(n2536), .CK(clk), .RN(rst_n), .Q(
        w_matrix[899]) );
  DFFRHQX1 w_matrix_reg_0__1__7_ ( .D(n2436), .CK(clk), .RN(rst_n), .Q(
        w_matrix[999]) );
  DFFRHQX1 w_matrix_reg_0__5__7_ ( .D(n2500), .CK(clk), .RN(rst_n), .Q(
        w_matrix[935]) );
  DFFRHQX1 w_matrix_reg_0__1__6_ ( .D(n2437), .CK(clk), .RN(rst_n), .Q(
        w_matrix[998]) );
  DFFRHQX1 w_matrix_reg_0__5__6_ ( .D(n2501), .CK(clk), .RN(rst_n), .Q(
        w_matrix[934]) );
  DFFRHQX1 w_matrix_reg_0__1__5_ ( .D(n2438), .CK(clk), .RN(rst_n), .Q(
        w_matrix[997]) );
  DFFRHQX1 w_matrix_reg_0__5__5_ ( .D(n2502), .CK(clk), .RN(rst_n), .Q(
        w_matrix[933]) );
  DFFRHQX1 w_matrix_reg_0__1__4_ ( .D(n2439), .CK(clk), .RN(rst_n), .Q(
        w_matrix[996]) );
  DFFRHQX1 w_matrix_reg_0__5__4_ ( .D(n2503), .CK(clk), .RN(rst_n), .Q(
        w_matrix[932]) );
  DFFRHQX1 w_matrix_reg_0__1__3_ ( .D(n2440), .CK(clk), .RN(rst_n), .Q(
        w_matrix[995]) );
  DFFRHQX1 w_matrix_reg_0__5__3_ ( .D(n2504), .CK(clk), .RN(rst_n), .Q(
        w_matrix[931]) );
  DFFRHQX1 w_matrix_reg_0__1__2_ ( .D(n2441), .CK(clk), .RN(rst_n), .Q(
        w_matrix[994]) );
  DFFRHQX1 w_matrix_reg_0__5__2_ ( .D(n2505), .CK(clk), .RN(rst_n), .Q(
        w_matrix[930]) );
  DFFRHQX1 w_matrix_reg_0__1__1_ ( .D(n2442), .CK(clk), .RN(rst_n), .Q(
        w_matrix[993]) );
  DFFRHQX1 w_matrix_reg_0__5__1_ ( .D(n2506), .CK(clk), .RN(rst_n), .Q(
        w_matrix[929]) );
  DFFRHQX1 w_matrix_reg_0__3__2_ ( .D(n2473), .CK(clk), .RN(rst_n), .Q(
        w_matrix[962]) );
  DFFRHQX1 w_matrix_reg_0__7__2_ ( .D(n2537), .CK(clk), .RN(rst_n), .Q(
        w_matrix[898]) );
  DFFRHQX1 w_matrix_reg_1__2__13_ ( .D(n2574), .CK(clk), .RN(rst_n), .Q(
        w_matrix[861]) );
  DFFRHQX1 w_matrix_reg_1__6__13_ ( .D(n2638), .CK(clk), .RN(rst_n), .Q(
        w_matrix[797]) );
  DFFRHQX1 w_matrix_reg_2__2__13_ ( .D(n2702), .CK(clk), .RN(rst_n), .Q(
        w_matrix[733]) );
  DFFRHQX1 w_matrix_reg_2__6__13_ ( .D(n2766), .CK(clk), .RN(rst_n), .Q(
        w_matrix[669]) );
  DFFRHQX1 w_matrix_reg_3__2__13_ ( .D(n2830), .CK(clk), .RN(rst_n), .Q(
        w_matrix[605]) );
  DFFRHQX1 w_matrix_reg_3__6__13_ ( .D(n2894), .CK(clk), .RN(rst_n), .Q(
        w_matrix[541]) );
  DFFRHQX1 w_matrix_reg_4__2__13_ ( .D(n2958), .CK(clk), .RN(rst_n), .Q(
        w_matrix[477]) );
  DFFRHQX1 w_matrix_reg_4__6__13_ ( .D(n3022), .CK(clk), .RN(rst_n), .Q(
        w_matrix[413]) );
  DFFRHQX1 w_matrix_reg_5__2__13_ ( .D(n3086), .CK(clk), .RN(rst_n), .Q(
        w_matrix[349]) );
  DFFRHQX1 w_matrix_reg_5__6__13_ ( .D(n3150), .CK(clk), .RN(rst_n), .Q(
        w_matrix[285]) );
  DFFRHQX1 w_matrix_reg_6__2__13_ ( .D(n3214), .CK(clk), .RN(rst_n), .Q(
        w_matrix[221]) );
  DFFRHQX1 w_matrix_reg_6__6__13_ ( .D(n3278), .CK(clk), .RN(rst_n), .Q(
        w_matrix[157]) );
  DFFRHQX1 w_matrix_reg_7__2__13_ ( .D(n3342), .CK(clk), .RN(rst_n), .Q(
        w_matrix[93]) );
  DFFRHQX1 w_matrix_reg_7__6__13_ ( .D(n3406), .CK(clk), .RN(rst_n), .Q(
        w_matrix[29]) );
  DFFRHQX1 w_matrix_reg_1__2__12_ ( .D(n2575), .CK(clk), .RN(rst_n), .Q(
        w_matrix[860]) );
  DFFRHQX1 w_matrix_reg_1__6__12_ ( .D(n2639), .CK(clk), .RN(rst_n), .Q(
        w_matrix[796]) );
  DFFRHQX1 w_matrix_reg_2__2__12_ ( .D(n2703), .CK(clk), .RN(rst_n), .Q(
        w_matrix[732]) );
  DFFRHQX1 w_matrix_reg_2__6__12_ ( .D(n2767), .CK(clk), .RN(rst_n), .Q(
        w_matrix[668]) );
  DFFRHQX1 w_matrix_reg_3__2__12_ ( .D(n2831), .CK(clk), .RN(rst_n), .Q(
        w_matrix[604]) );
  DFFRHQX1 w_matrix_reg_3__6__12_ ( .D(n2895), .CK(clk), .RN(rst_n), .Q(
        w_matrix[540]) );
  DFFRHQX1 w_matrix_reg_4__2__12_ ( .D(n2959), .CK(clk), .RN(rst_n), .Q(
        w_matrix[476]) );
  DFFRHQX1 w_matrix_reg_4__6__12_ ( .D(n3023), .CK(clk), .RN(rst_n), .Q(
        w_matrix[412]) );
  DFFRHQX1 w_matrix_reg_5__2__12_ ( .D(n3087), .CK(clk), .RN(rst_n), .Q(
        w_matrix[348]) );
  DFFRHQX1 w_matrix_reg_5__6__12_ ( .D(n3151), .CK(clk), .RN(rst_n), .Q(
        w_matrix[284]) );
  DFFRHQX1 w_matrix_reg_6__2__12_ ( .D(n3215), .CK(clk), .RN(rst_n), .Q(
        w_matrix[220]) );
  DFFRHQX1 w_matrix_reg_6__6__12_ ( .D(n3279), .CK(clk), .RN(rst_n), .Q(
        w_matrix[156]) );
  DFFRHQX1 w_matrix_reg_7__2__12_ ( .D(n3343), .CK(clk), .RN(rst_n), .Q(
        w_matrix[92]) );
  DFFRHQX1 w_matrix_reg_7__6__12_ ( .D(n3407), .CK(clk), .RN(rst_n), .Q(
        w_matrix[28]) );
  DFFRHQX1 w_matrix_reg_1__2__11_ ( .D(n2576), .CK(clk), .RN(rst_n), .Q(
        w_matrix[859]) );
  DFFRHQX1 w_matrix_reg_1__6__11_ ( .D(n2640), .CK(clk), .RN(rst_n), .Q(
        w_matrix[795]) );
  DFFRHQX1 w_matrix_reg_2__2__11_ ( .D(n2704), .CK(clk), .RN(rst_n), .Q(
        w_matrix[731]) );
  DFFRHQX1 w_matrix_reg_2__6__11_ ( .D(n2768), .CK(clk), .RN(rst_n), .Q(
        w_matrix[667]) );
  DFFRHQX1 w_matrix_reg_3__2__11_ ( .D(n2832), .CK(clk), .RN(rst_n), .Q(
        w_matrix[603]) );
  DFFRHQX1 w_matrix_reg_3__6__11_ ( .D(n2896), .CK(clk), .RN(rst_n), .Q(
        w_matrix[539]) );
  DFFRHQX1 w_matrix_reg_4__2__11_ ( .D(n2960), .CK(clk), .RN(rst_n), .Q(
        w_matrix[475]) );
  DFFRHQX1 w_matrix_reg_4__6__11_ ( .D(n3024), .CK(clk), .RN(rst_n), .Q(
        w_matrix[411]) );
  DFFRHQX1 w_matrix_reg_5__2__11_ ( .D(n3088), .CK(clk), .RN(rst_n), .Q(
        w_matrix[347]) );
  DFFRHQX1 w_matrix_reg_5__6__11_ ( .D(n3152), .CK(clk), .RN(rst_n), .Q(
        w_matrix[283]) );
  DFFRHQX1 w_matrix_reg_6__2__11_ ( .D(n3216), .CK(clk), .RN(rst_n), .Q(
        w_matrix[219]) );
  DFFRHQX1 w_matrix_reg_6__6__11_ ( .D(n3280), .CK(clk), .RN(rst_n), .Q(
        w_matrix[155]) );
  DFFRHQX1 w_matrix_reg_7__2__11_ ( .D(n3344), .CK(clk), .RN(rst_n), .Q(
        w_matrix[91]) );
  DFFRHQX1 w_matrix_reg_7__6__11_ ( .D(n3408), .CK(clk), .RN(rst_n), .Q(
        w_matrix[27]) );
  DFFRHQX1 w_matrix_reg_0__2__7_ ( .D(n2452), .CK(clk), .RN(rst_n), .Q(
        w_matrix[983]) );
  DFFRHQX1 w_matrix_reg_0__6__7_ ( .D(n2516), .CK(clk), .RN(rst_n), .Q(
        w_matrix[919]) );
  DFFRHQX1 w_matrix_reg_0__2__6_ ( .D(n2453), .CK(clk), .RN(rst_n), .Q(
        w_matrix[982]) );
  DFFRHQX1 w_matrix_reg_0__6__6_ ( .D(n2517), .CK(clk), .RN(rst_n), .Q(
        w_matrix[918]) );
  DFFRHQX1 w_matrix_reg_0__2__5_ ( .D(n2454), .CK(clk), .RN(rst_n), .Q(
        w_matrix[981]) );
  DFFRHQX1 w_matrix_reg_0__6__5_ ( .D(n2518), .CK(clk), .RN(rst_n), .Q(
        w_matrix[917]) );
  DFFRHQX1 w_matrix_reg_0__2__4_ ( .D(n2455), .CK(clk), .RN(rst_n), .Q(
        w_matrix[980]) );
  DFFRHQX1 w_matrix_reg_0__6__4_ ( .D(n2519), .CK(clk), .RN(rst_n), .Q(
        w_matrix[916]) );
  DFFRHQX1 w_matrix_reg_0__3__1_ ( .D(n2474), .CK(clk), .RN(rst_n), .Q(
        w_matrix[961]) );
  DFFRHQX1 w_matrix_reg_0__7__1_ ( .D(n2538), .CK(clk), .RN(rst_n), .Q(
        w_matrix[897]) );
  DFFRHQX1 w_matrix_reg_0__2__3_ ( .D(n2456), .CK(clk), .RN(rst_n), .Q(
        w_matrix[979]) );
  DFFRHQX1 w_matrix_reg_0__6__3_ ( .D(n2520), .CK(clk), .RN(rst_n), .Q(
        w_matrix[915]) );
  DFFRHQX1 w_matrix_reg_0__2__2_ ( .D(n2457), .CK(clk), .RN(rst_n), .Q(
        w_matrix[978]) );
  DFFRHQX1 w_matrix_reg_0__6__2_ ( .D(n2521), .CK(clk), .RN(rst_n), .Q(
        w_matrix[914]) );
  DFFRHQX1 w_matrix_reg_0__2__1_ ( .D(n2458), .CK(clk), .RN(rst_n), .Q(
        w_matrix[977]) );
  DFFRHQX1 w_matrix_reg_0__6__1_ ( .D(n2522), .CK(clk), .RN(rst_n), .Q(
        w_matrix[913]) );
  DFFRHQX1 w_matrix_reg_1__3__13_ ( .D(n2590), .CK(clk), .RN(rst_n), .Q(
        w_matrix[845]) );
  DFFRHQX1 w_matrix_reg_1__7__13_ ( .D(n2654), .CK(clk), .RN(rst_n), .Q(
        w_matrix[781]) );
  DFFRHQX1 w_matrix_reg_2__3__13_ ( .D(n2718), .CK(clk), .RN(rst_n), .Q(
        w_matrix[717]) );
  DFFRHQX1 w_matrix_reg_2__7__13_ ( .D(n2782), .CK(clk), .RN(rst_n), .Q(
        w_matrix[653]) );
  DFFRHQX1 w_matrix_reg_3__3__13_ ( .D(n2846), .CK(clk), .RN(rst_n), .Q(
        w_matrix[589]) );
  DFFRHQX1 w_matrix_reg_3__7__13_ ( .D(n2910), .CK(clk), .RN(rst_n), .Q(
        w_matrix[525]) );
  DFFRHQX1 w_matrix_reg_4__3__13_ ( .D(n2974), .CK(clk), .RN(rst_n), .Q(
        w_matrix[461]) );
  DFFRHQX1 w_matrix_reg_4__7__13_ ( .D(n3038), .CK(clk), .RN(rst_n), .Q(
        w_matrix[397]) );
  DFFRHQX1 w_matrix_reg_5__3__13_ ( .D(n3102), .CK(clk), .RN(rst_n), .Q(
        w_matrix[333]) );
  DFFRHQX1 w_matrix_reg_5__7__13_ ( .D(n3166), .CK(clk), .RN(rst_n), .Q(
        w_matrix[269]) );
  DFFRHQX1 w_matrix_reg_6__3__13_ ( .D(n3230), .CK(clk), .RN(rst_n), .Q(
        w_matrix[205]) );
  DFFRHQX1 w_matrix_reg_6__7__13_ ( .D(n3294), .CK(clk), .RN(rst_n), .Q(
        w_matrix[141]) );
  DFFRHQX1 w_matrix_reg_7__3__13_ ( .D(n3358), .CK(clk), .RN(rst_n), .Q(
        w_matrix[77]) );
  DFFRHQX1 w_matrix_reg_7__7__13_ ( .D(n3422), .CK(clk), .RN(rst_n), .Q(
        w_matrix[13]) );
  DFFRHQX1 w_matrix_reg_1__3__12_ ( .D(n2591), .CK(clk), .RN(rst_n), .Q(
        w_matrix[844]) );
  DFFRHQX1 w_matrix_reg_1__7__12_ ( .D(n2655), .CK(clk), .RN(rst_n), .Q(
        w_matrix[780]) );
  DFFRHQX1 w_matrix_reg_2__3__12_ ( .D(n2719), .CK(clk), .RN(rst_n), .Q(
        w_matrix[716]) );
  DFFRHQX1 w_matrix_reg_2__7__12_ ( .D(n2783), .CK(clk), .RN(rst_n), .Q(
        w_matrix[652]) );
  DFFRHQX1 w_matrix_reg_3__3__12_ ( .D(n2847), .CK(clk), .RN(rst_n), .Q(
        w_matrix[588]) );
  DFFRHQX1 w_matrix_reg_3__7__12_ ( .D(n2911), .CK(clk), .RN(rst_n), .Q(
        w_matrix[524]) );
  DFFRHQX1 w_matrix_reg_4__3__12_ ( .D(n2975), .CK(clk), .RN(rst_n), .Q(
        w_matrix[460]) );
  DFFRHQX1 w_matrix_reg_4__7__12_ ( .D(n3039), .CK(clk), .RN(rst_n), .Q(
        w_matrix[396]) );
  DFFRHQX1 w_matrix_reg_5__3__12_ ( .D(n3103), .CK(clk), .RN(rst_n), .Q(
        w_matrix[332]) );
  DFFRHQX1 w_matrix_reg_5__7__12_ ( .D(n3167), .CK(clk), .RN(rst_n), .Q(
        w_matrix[268]) );
  DFFRHQX1 w_matrix_reg_6__3__12_ ( .D(n3231), .CK(clk), .RN(rst_n), .Q(
        w_matrix[204]) );
  DFFRHQX1 w_matrix_reg_6__7__12_ ( .D(n3295), .CK(clk), .RN(rst_n), .Q(
        w_matrix[140]) );
  DFFRHQX1 w_matrix_reg_7__3__12_ ( .D(n3359), .CK(clk), .RN(rst_n), .Q(
        w_matrix[76]) );
  DFFRHQX1 w_matrix_reg_7__7__12_ ( .D(n3423), .CK(clk), .RN(rst_n), .Q(
        w_matrix[12]) );
  DFFRHQX1 w_matrix_reg_1__3__11_ ( .D(n2592), .CK(clk), .RN(rst_n), .Q(
        w_matrix[843]) );
  DFFRHQX1 w_matrix_reg_1__7__11_ ( .D(n2656), .CK(clk), .RN(rst_n), .Q(
        w_matrix[779]) );
  DFFRHQX1 w_matrix_reg_2__3__11_ ( .D(n2720), .CK(clk), .RN(rst_n), .Q(
        w_matrix[715]) );
  DFFRHQX1 w_matrix_reg_2__7__11_ ( .D(n2784), .CK(clk), .RN(rst_n), .Q(
        w_matrix[651]) );
  DFFRHQX1 w_matrix_reg_3__3__11_ ( .D(n2848), .CK(clk), .RN(rst_n), .Q(
        w_matrix[587]) );
  DFFRHQX1 w_matrix_reg_3__7__11_ ( .D(n2912), .CK(clk), .RN(rst_n), .Q(
        w_matrix[523]) );
  DFFRHQX1 w_matrix_reg_4__3__11_ ( .D(n2976), .CK(clk), .RN(rst_n), .Q(
        w_matrix[459]) );
  DFFRHQX1 w_matrix_reg_4__7__11_ ( .D(n3040), .CK(clk), .RN(rst_n), .Q(
        w_matrix[395]) );
  DFFRHQX1 w_matrix_reg_5__3__11_ ( .D(n3104), .CK(clk), .RN(rst_n), .Q(
        w_matrix[331]) );
  DFFRHQX1 w_matrix_reg_5__7__11_ ( .D(n3168), .CK(clk), .RN(rst_n), .Q(
        w_matrix[267]) );
  DFFRHQX1 w_matrix_reg_6__3__11_ ( .D(n3232), .CK(clk), .RN(rst_n), .Q(
        w_matrix[203]) );
  DFFRHQX1 w_matrix_reg_6__7__11_ ( .D(n3296), .CK(clk), .RN(rst_n), .Q(
        w_matrix[139]) );
  DFFRHQX1 w_matrix_reg_7__3__11_ ( .D(n3360), .CK(clk), .RN(rst_n), .Q(
        w_matrix[75]) );
  DFFRHQX1 w_matrix_reg_7__7__11_ ( .D(n3424), .CK(clk), .RN(rst_n), .Q(
        w_matrix[11]) );
  DFFRHQX1 inA11_reg_0_ ( .D(N11394), .CK(clk), .RN(rst_n), .Q(inA11[0]) );
  DFFRHQX1 w_matrix_reg_1__0__14_ ( .D(n2541), .CK(clk), .RN(rst_n), .Q(
        w_matrix[894]) );
  DFFRX1 w_matrix_reg_1__1__9_ ( .D(n2562), .CK(clk), .RN(rst_n), .Q(
        w_matrix[873]), .QN(n664) );
  DFFRX1 w_matrix_reg_1__1__8_ ( .D(n2563), .CK(clk), .RN(rst_n), .Q(
        w_matrix[872]), .QN(n665) );
  DFFRX1 w_matrix_reg_1__1__12_ ( .D(n2559), .CK(clk), .RN(rst_n), .Q(
        w_matrix[876]), .QN(n661) );
  DFFRX1 w_matrix_reg_1__1__11_ ( .D(n2560), .CK(clk), .RN(rst_n), .Q(
        w_matrix[875]), .QN(n662) );
  DFFRX1 w_matrix_reg_1__1__10_ ( .D(n2561), .CK(clk), .RN(rst_n), .Q(
        w_matrix[874]), .QN(n663) );
  DFFRHQX1 inA41_reg_8_ ( .D(N11689), .CK(clk), .RN(rst_n), .Q(inA41[8]) );
  DFFRHQX1 inA81_reg_8_ ( .D(N12068), .CK(clk), .RN(rst_n), .Q(inA81[8]) );
  DFFRHQX1 inA51_reg_10_ ( .D(N11783), .CK(clk), .RN(rst_n), .Q(inA51[10]) );
  DFFRHQX1 inA51_reg_8_ ( .D(N11781), .CK(clk), .RN(rst_n), .Q(inA51[8]) );
  DFFRHQX1 inA61_reg_10_ ( .D(N11880), .CK(clk), .RN(rst_n), .Q(inA61[10]) );
  DFFRHQX1 inA21_reg_8_ ( .D(N11498), .CK(clk), .RN(rst_n), .Q(inA21[8]) );
  DFFRHQX1 inA61_reg_8_ ( .D(N11878), .CK(clk), .RN(rst_n), .Q(inA61[8]) );
  DFFRHQX1 inA31_reg_10_ ( .D(N11594), .CK(clk), .RN(rst_n), .Q(inA31[10]) );
  DFFRHQX1 inA71_reg_10_ ( .D(N11974), .CK(clk), .RN(rst_n), .Q(inA71[10]) );
  DFFRHQX1 inA31_reg_8_ ( .D(N11592), .CK(clk), .RN(rst_n), .Q(inA31[8]) );
  DFFRHQX1 inA71_reg_8_ ( .D(N11972), .CK(clk), .RN(rst_n), .Q(inA71[8]) );
  DFFRHQX1 inA21_reg_10_ ( .D(N11500), .CK(clk), .RN(rst_n), .Q(inA21[10]) );
  DFFRHQX1 inA41_reg_10_ ( .D(N11691), .CK(clk), .RN(rst_n), .Q(inA41[10]) );
  DFFRHQX1 inA81_reg_10_ ( .D(N12070), .CK(clk), .RN(rst_n), .Q(inA81[10]) );
  DFFRHQX1 inA41_reg_9_ ( .D(N11690), .CK(clk), .RN(rst_n), .Q(inA41[9]) );
  DFFRHQX1 inA81_reg_9_ ( .D(N12069), .CK(clk), .RN(rst_n), .Q(inA81[9]) );
  DFFRHQX1 inA51_reg_13_ ( .D(N11786), .CK(clk), .RN(rst_n), .Q(inA51[13]) );
  DFFRHQX1 inA51_reg_11_ ( .D(N11784), .CK(clk), .RN(rst_n), .Q(inA51[11]) );
  DFFRHQX1 inA51_reg_9_ ( .D(N11782), .CK(clk), .RN(rst_n), .Q(inA51[9]) );
  DFFRHQX1 inA61_reg_13_ ( .D(N11883), .CK(clk), .RN(rst_n), .Q(inA61[13]) );
  DFFRHQX1 inA61_reg_11_ ( .D(N11881), .CK(clk), .RN(rst_n), .Q(inA61[11]) );
  DFFRHQX1 inA21_reg_9_ ( .D(N11499), .CK(clk), .RN(rst_n), .Q(inA21[9]) );
  DFFRHQX1 inA61_reg_9_ ( .D(N11879), .CK(clk), .RN(rst_n), .Q(inA61[9]) );
  DFFRHQX1 inA31_reg_13_ ( .D(N11597), .CK(clk), .RN(rst_n), .Q(inA31[13]) );
  DFFRHQX1 inA71_reg_13_ ( .D(N11977), .CK(clk), .RN(rst_n), .Q(inA71[13]) );
  DFFRHQX1 inA31_reg_11_ ( .D(N11595), .CK(clk), .RN(rst_n), .Q(inA31[11]) );
  DFFRHQX1 inA71_reg_11_ ( .D(N11975), .CK(clk), .RN(rst_n), .Q(inA71[11]) );
  DFFRHQX1 inA31_reg_9_ ( .D(N11593), .CK(clk), .RN(rst_n), .Q(inA31[9]) );
  DFFRHQX1 inA71_reg_9_ ( .D(N11973), .CK(clk), .RN(rst_n), .Q(inA71[9]) );
  DFFRHQX1 inA11_reg_3_ ( .D(N11397), .CK(clk), .RN(rst_n), .Q(inA11[3]) );
  DFFRHQX1 inA11_reg_1_ ( .D(N11395), .CK(clk), .RN(rst_n), .Q(inA11[1]) );
  DFFRHQX1 inA21_reg_13_ ( .D(N11503), .CK(clk), .RN(rst_n), .Q(inA21[13]) );
  DFFRHQX1 inA41_reg_13_ ( .D(N11694), .CK(clk), .RN(rst_n), .Q(inA41[13]) );
  DFFRHQX1 inA81_reg_13_ ( .D(N12073), .CK(clk), .RN(rst_n), .Q(inA81[13]) );
  DFFRHQX1 inA21_reg_11_ ( .D(N11501), .CK(clk), .RN(rst_n), .Q(inA21[11]) );
  DFFRHQX1 inA41_reg_11_ ( .D(N11692), .CK(clk), .RN(rst_n), .Q(inA41[11]) );
  DFFRHQX1 inA81_reg_11_ ( .D(N12071), .CK(clk), .RN(rst_n), .Q(inA81[11]) );
  DFFRHQX1 w_matrix_reg_1__3__9_ ( .D(n2594), .CK(clk), .RN(rst_n), .Q(
        w_matrix[841]) );
  DFFRHQX1 w_matrix_reg_1__7__9_ ( .D(n2658), .CK(clk), .RN(rst_n), .Q(
        w_matrix[777]) );
  DFFRHQX1 w_matrix_reg_2__3__9_ ( .D(n2722), .CK(clk), .RN(rst_n), .Q(
        w_matrix[713]) );
  DFFRHQX1 w_matrix_reg_2__7__9_ ( .D(n2786), .CK(clk), .RN(rst_n), .Q(
        w_matrix[649]) );
  DFFRHQX1 w_matrix_reg_3__3__9_ ( .D(n2850), .CK(clk), .RN(rst_n), .Q(
        w_matrix[585]) );
  DFFRHQX1 w_matrix_reg_3__7__9_ ( .D(n2914), .CK(clk), .RN(rst_n), .Q(
        w_matrix[521]) );
  DFFRHQX1 w_matrix_reg_4__3__9_ ( .D(n2978), .CK(clk), .RN(rst_n), .Q(
        w_matrix[457]) );
  DFFRHQX1 w_matrix_reg_4__7__9_ ( .D(n3042), .CK(clk), .RN(rst_n), .Q(
        w_matrix[393]) );
  DFFRHQX1 w_matrix_reg_5__3__9_ ( .D(n3106), .CK(clk), .RN(rst_n), .Q(
        w_matrix[329]) );
  DFFRHQX1 w_matrix_reg_5__7__9_ ( .D(n3170), .CK(clk), .RN(rst_n), .Q(
        w_matrix[265]) );
  DFFRHQX1 w_matrix_reg_6__3__9_ ( .D(n3234), .CK(clk), .RN(rst_n), .Q(
        w_matrix[201]) );
  DFFRHQX1 w_matrix_reg_6__7__9_ ( .D(n3298), .CK(clk), .RN(rst_n), .Q(
        w_matrix[137]) );
  DFFRHQX1 w_matrix_reg_7__3__9_ ( .D(n3362), .CK(clk), .RN(rst_n), .Q(
        w_matrix[73]) );
  DFFRHQX1 w_matrix_reg_7__7__9_ ( .D(n3426), .CK(clk), .RN(rst_n), .Q(
        w_matrix[9]) );
  DFFRHQX1 w_matrix_reg_1__3__8_ ( .D(n2595), .CK(clk), .RN(rst_n), .Q(
        w_matrix[840]) );
  DFFRHQX1 w_matrix_reg_1__7__8_ ( .D(n2659), .CK(clk), .RN(rst_n), .Q(
        w_matrix[776]) );
  DFFRHQX1 w_matrix_reg_2__3__8_ ( .D(n2723), .CK(clk), .RN(rst_n), .Q(
        w_matrix[712]) );
  DFFRHQX1 w_matrix_reg_2__7__8_ ( .D(n2787), .CK(clk), .RN(rst_n), .Q(
        w_matrix[648]) );
  DFFRHQX1 w_matrix_reg_3__3__8_ ( .D(n2851), .CK(clk), .RN(rst_n), .Q(
        w_matrix[584]) );
  DFFRHQX1 w_matrix_reg_3__7__8_ ( .D(n2915), .CK(clk), .RN(rst_n), .Q(
        w_matrix[520]) );
  DFFRHQX1 w_matrix_reg_4__3__8_ ( .D(n2979), .CK(clk), .RN(rst_n), .Q(
        w_matrix[456]) );
  DFFRHQX1 w_matrix_reg_4__7__8_ ( .D(n3043), .CK(clk), .RN(rst_n), .Q(
        w_matrix[392]) );
  DFFRHQX1 w_matrix_reg_5__3__8_ ( .D(n3107), .CK(clk), .RN(rst_n), .Q(
        w_matrix[328]) );
  DFFRHQX1 w_matrix_reg_5__7__8_ ( .D(n3171), .CK(clk), .RN(rst_n), .Q(
        w_matrix[264]) );
  DFFRHQX1 w_matrix_reg_6__3__8_ ( .D(n3235), .CK(clk), .RN(rst_n), .Q(
        w_matrix[200]) );
  DFFRHQX1 w_matrix_reg_6__7__8_ ( .D(n3299), .CK(clk), .RN(rst_n), .Q(
        w_matrix[136]) );
  DFFRHQX1 w_matrix_reg_7__3__8_ ( .D(n3363), .CK(clk), .RN(rst_n), .Q(
        w_matrix[72]) );
  DFFRHQX1 w_matrix_reg_7__7__8_ ( .D(n3427), .CK(clk), .RN(rst_n), .Q(
        w_matrix[8]) );
  DFFRHQX1 w_matrix_reg_1__4__10_ ( .D(n2609), .CK(clk), .RN(rst_n), .Q(
        w_matrix[826]) );
  DFFRHQX1 w_matrix_reg_2__0__10_ ( .D(n2673), .CK(clk), .RN(rst_n), .Q(
        w_matrix[762]) );
  DFFRHQX1 w_matrix_reg_2__4__10_ ( .D(n2737), .CK(clk), .RN(rst_n), .Q(
        w_matrix[698]) );
  DFFRHQX1 w_matrix_reg_3__0__10_ ( .D(n2801), .CK(clk), .RN(rst_n), .Q(
        w_matrix[634]) );
  DFFRHQX1 w_matrix_reg_3__4__10_ ( .D(n2865), .CK(clk), .RN(rst_n), .Q(
        w_matrix[570]) );
  DFFRHQX1 w_matrix_reg_4__0__10_ ( .D(n2929), .CK(clk), .RN(rst_n), .Q(
        w_matrix[506]) );
  DFFRHQX1 w_matrix_reg_4__4__10_ ( .D(n2993), .CK(clk), .RN(rst_n), .Q(
        w_matrix[442]) );
  DFFRHQX1 w_matrix_reg_5__0__10_ ( .D(n3057), .CK(clk), .RN(rst_n), .Q(
        w_matrix[378]) );
  DFFRHQX1 w_matrix_reg_5__4__10_ ( .D(n3121), .CK(clk), .RN(rst_n), .Q(
        w_matrix[314]) );
  DFFRHQX1 w_matrix_reg_6__0__10_ ( .D(n3185), .CK(clk), .RN(rst_n), .Q(
        w_matrix[250]) );
  DFFRHQX1 w_matrix_reg_6__4__10_ ( .D(n3249), .CK(clk), .RN(rst_n), .Q(
        w_matrix[186]) );
  DFFRHQX1 w_matrix_reg_7__0__10_ ( .D(n3313), .CK(clk), .RN(rst_n), .Q(
        w_matrix[122]) );
  DFFRHQX1 w_matrix_reg_7__4__10_ ( .D(n3377), .CK(clk), .RN(rst_n), .Q(
        w_matrix[58]) );
  DFFRHQX1 w_matrix_reg_1__4__9_ ( .D(n2610), .CK(clk), .RN(rst_n), .Q(
        w_matrix[825]) );
  DFFRHQX1 w_matrix_reg_2__0__9_ ( .D(n2674), .CK(clk), .RN(rst_n), .Q(
        w_matrix[761]) );
  DFFRHQX1 w_matrix_reg_2__4__9_ ( .D(n2738), .CK(clk), .RN(rst_n), .Q(
        w_matrix[697]) );
  DFFRHQX1 w_matrix_reg_3__0__9_ ( .D(n2802), .CK(clk), .RN(rst_n), .Q(
        w_matrix[633]) );
  DFFRHQX1 w_matrix_reg_3__4__9_ ( .D(n2866), .CK(clk), .RN(rst_n), .Q(
        w_matrix[569]) );
  DFFRHQX1 w_matrix_reg_4__0__9_ ( .D(n2930), .CK(clk), .RN(rst_n), .Q(
        w_matrix[505]) );
  DFFRHQX1 w_matrix_reg_4__4__9_ ( .D(n2994), .CK(clk), .RN(rst_n), .Q(
        w_matrix[441]) );
  DFFRHQX1 w_matrix_reg_5__0__9_ ( .D(n3058), .CK(clk), .RN(rst_n), .Q(
        w_matrix[377]) );
  DFFRHQX1 w_matrix_reg_5__4__9_ ( .D(n3122), .CK(clk), .RN(rst_n), .Q(
        w_matrix[313]) );
  DFFRHQX1 w_matrix_reg_6__0__9_ ( .D(n3186), .CK(clk), .RN(rst_n), .Q(
        w_matrix[249]) );
  DFFRHQX1 w_matrix_reg_6__4__9_ ( .D(n3250), .CK(clk), .RN(rst_n), .Q(
        w_matrix[185]) );
  DFFRHQX1 w_matrix_reg_7__0__9_ ( .D(n3314), .CK(clk), .RN(rst_n), .Q(
        w_matrix[121]) );
  DFFRHQX1 w_matrix_reg_7__4__9_ ( .D(n3378), .CK(clk), .RN(rst_n), .Q(
        w_matrix[57]) );
  DFFRHQX1 w_matrix_reg_1__4__8_ ( .D(n2611), .CK(clk), .RN(rst_n), .Q(
        w_matrix[824]) );
  DFFRHQX1 w_matrix_reg_2__0__8_ ( .D(n2675), .CK(clk), .RN(rst_n), .Q(
        w_matrix[760]) );
  DFFRHQX1 w_matrix_reg_2__4__8_ ( .D(n2739), .CK(clk), .RN(rst_n), .Q(
        w_matrix[696]) );
  DFFRHQX1 w_matrix_reg_3__0__8_ ( .D(n2803), .CK(clk), .RN(rst_n), .Q(
        w_matrix[632]) );
  DFFRHQX1 w_matrix_reg_3__4__8_ ( .D(n2867), .CK(clk), .RN(rst_n), .Q(
        w_matrix[568]) );
  DFFRHQX1 w_matrix_reg_4__0__8_ ( .D(n2931), .CK(clk), .RN(rst_n), .Q(
        w_matrix[504]) );
  DFFRHQX1 w_matrix_reg_4__4__8_ ( .D(n2995), .CK(clk), .RN(rst_n), .Q(
        w_matrix[440]) );
  DFFRHQX1 w_matrix_reg_5__0__8_ ( .D(n3059), .CK(clk), .RN(rst_n), .Q(
        w_matrix[376]) );
  DFFRHQX1 w_matrix_reg_5__4__8_ ( .D(n3123), .CK(clk), .RN(rst_n), .Q(
        w_matrix[312]) );
  DFFRHQX1 w_matrix_reg_6__0__8_ ( .D(n3187), .CK(clk), .RN(rst_n), .Q(
        w_matrix[248]) );
  DFFRHQX1 w_matrix_reg_6__4__8_ ( .D(n3251), .CK(clk), .RN(rst_n), .Q(
        w_matrix[184]) );
  DFFRHQX1 w_matrix_reg_7__0__8_ ( .D(n3315), .CK(clk), .RN(rst_n), .Q(
        w_matrix[120]) );
  DFFRHQX1 w_matrix_reg_7__4__8_ ( .D(n3379), .CK(clk), .RN(rst_n), .Q(
        w_matrix[56]) );
  DFFRHQX1 w_matrix_reg_1__5__10_ ( .D(n2625), .CK(clk), .RN(rst_n), .Q(
        w_matrix[810]) );
  DFFRHQX1 w_matrix_reg_2__1__10_ ( .D(n2689), .CK(clk), .RN(rst_n), .Q(
        w_matrix[746]) );
  DFFRHQX1 w_matrix_reg_2__5__10_ ( .D(n2753), .CK(clk), .RN(rst_n), .Q(
        w_matrix[682]) );
  DFFRHQX1 w_matrix_reg_3__1__10_ ( .D(n2817), .CK(clk), .RN(rst_n), .Q(
        w_matrix[618]) );
  DFFRHQX1 w_matrix_reg_3__5__10_ ( .D(n2881), .CK(clk), .RN(rst_n), .Q(
        w_matrix[554]) );
  DFFRHQX1 w_matrix_reg_4__1__10_ ( .D(n2945), .CK(clk), .RN(rst_n), .Q(
        w_matrix[490]) );
  DFFRHQX1 w_matrix_reg_4__5__10_ ( .D(n3009), .CK(clk), .RN(rst_n), .Q(
        w_matrix[426]) );
  DFFRHQX1 w_matrix_reg_5__1__10_ ( .D(n3073), .CK(clk), .RN(rst_n), .Q(
        w_matrix[362]) );
  DFFRHQX1 w_matrix_reg_5__5__10_ ( .D(n3137), .CK(clk), .RN(rst_n), .Q(
        w_matrix[298]) );
  DFFRHQX1 w_matrix_reg_6__1__10_ ( .D(n3201), .CK(clk), .RN(rst_n), .Q(
        w_matrix[234]) );
  DFFRHQX1 w_matrix_reg_6__5__10_ ( .D(n3265), .CK(clk), .RN(rst_n), .Q(
        w_matrix[170]) );
  DFFRHQX1 w_matrix_reg_7__1__10_ ( .D(n3329), .CK(clk), .RN(rst_n), .Q(
        w_matrix[106]) );
  DFFRHQX1 w_matrix_reg_7__5__10_ ( .D(n3393), .CK(clk), .RN(rst_n), .Q(
        w_matrix[42]) );
  DFFRHQX1 w_matrix_reg_1__5__9_ ( .D(n2626), .CK(clk), .RN(rst_n), .Q(
        w_matrix[809]) );
  DFFRHQX1 w_matrix_reg_2__1__9_ ( .D(n2690), .CK(clk), .RN(rst_n), .Q(
        w_matrix[745]) );
  DFFRHQX1 w_matrix_reg_2__5__9_ ( .D(n2754), .CK(clk), .RN(rst_n), .Q(
        w_matrix[681]) );
  DFFRHQX1 w_matrix_reg_3__1__9_ ( .D(n2818), .CK(clk), .RN(rst_n), .Q(
        w_matrix[617]) );
  DFFRHQX1 w_matrix_reg_3__5__9_ ( .D(n2882), .CK(clk), .RN(rst_n), .Q(
        w_matrix[553]) );
  DFFRHQX1 w_matrix_reg_4__1__9_ ( .D(n2946), .CK(clk), .RN(rst_n), .Q(
        w_matrix[489]) );
  DFFRHQX1 w_matrix_reg_4__5__9_ ( .D(n3010), .CK(clk), .RN(rst_n), .Q(
        w_matrix[425]) );
  DFFRHQX1 w_matrix_reg_5__1__9_ ( .D(n3074), .CK(clk), .RN(rst_n), .Q(
        w_matrix[361]) );
  DFFRHQX1 w_matrix_reg_5__5__9_ ( .D(n3138), .CK(clk), .RN(rst_n), .Q(
        w_matrix[297]) );
  DFFRHQX1 w_matrix_reg_6__1__9_ ( .D(n3202), .CK(clk), .RN(rst_n), .Q(
        w_matrix[233]) );
  DFFRHQX1 w_matrix_reg_6__5__9_ ( .D(n3266), .CK(clk), .RN(rst_n), .Q(
        w_matrix[169]) );
  DFFRHQX1 w_matrix_reg_7__1__9_ ( .D(n3330), .CK(clk), .RN(rst_n), .Q(
        w_matrix[105]) );
  DFFRHQX1 w_matrix_reg_7__5__9_ ( .D(n3394), .CK(clk), .RN(rst_n), .Q(
        w_matrix[41]) );
  DFFRHQX1 w_matrix_reg_1__5__8_ ( .D(n2627), .CK(clk), .RN(rst_n), .Q(
        w_matrix[808]) );
  DFFRHQX1 w_matrix_reg_2__1__8_ ( .D(n2691), .CK(clk), .RN(rst_n), .Q(
        w_matrix[744]) );
  DFFRHQX1 w_matrix_reg_2__5__8_ ( .D(n2755), .CK(clk), .RN(rst_n), .Q(
        w_matrix[680]) );
  DFFRHQX1 w_matrix_reg_3__1__8_ ( .D(n2819), .CK(clk), .RN(rst_n), .Q(
        w_matrix[616]) );
  DFFRHQX1 w_matrix_reg_3__5__8_ ( .D(n2883), .CK(clk), .RN(rst_n), .Q(
        w_matrix[552]) );
  DFFRHQX1 w_matrix_reg_4__1__8_ ( .D(n2947), .CK(clk), .RN(rst_n), .Q(
        w_matrix[488]) );
  DFFRHQX1 w_matrix_reg_4__5__8_ ( .D(n3011), .CK(clk), .RN(rst_n), .Q(
        w_matrix[424]) );
  DFFRHQX1 w_matrix_reg_5__1__8_ ( .D(n3075), .CK(clk), .RN(rst_n), .Q(
        w_matrix[360]) );
  DFFRHQX1 w_matrix_reg_5__5__8_ ( .D(n3139), .CK(clk), .RN(rst_n), .Q(
        w_matrix[296]) );
  DFFRHQX1 w_matrix_reg_6__1__8_ ( .D(n3203), .CK(clk), .RN(rst_n), .Q(
        w_matrix[232]) );
  DFFRHQX1 w_matrix_reg_6__5__8_ ( .D(n3267), .CK(clk), .RN(rst_n), .Q(
        w_matrix[168]) );
  DFFRHQX1 w_matrix_reg_7__1__8_ ( .D(n3331), .CK(clk), .RN(rst_n), .Q(
        w_matrix[104]) );
  DFFRHQX1 w_matrix_reg_7__5__8_ ( .D(n3395), .CK(clk), .RN(rst_n), .Q(
        w_matrix[40]) );
  DFFRHQX1 w_matrix_reg_1__2__10_ ( .D(n2577), .CK(clk), .RN(rst_n), .Q(
        w_matrix[858]) );
  DFFRHQX1 w_matrix_reg_1__6__10_ ( .D(n2641), .CK(clk), .RN(rst_n), .Q(
        w_matrix[794]) );
  DFFRHQX1 w_matrix_reg_2__2__10_ ( .D(n2705), .CK(clk), .RN(rst_n), .Q(
        w_matrix[730]) );
  DFFRHQX1 w_matrix_reg_2__6__10_ ( .D(n2769), .CK(clk), .RN(rst_n), .Q(
        w_matrix[666]) );
  DFFRHQX1 w_matrix_reg_3__2__10_ ( .D(n2833), .CK(clk), .RN(rst_n), .Q(
        w_matrix[602]) );
  DFFRHQX1 w_matrix_reg_3__6__10_ ( .D(n2897), .CK(clk), .RN(rst_n), .Q(
        w_matrix[538]) );
  DFFRHQX1 w_matrix_reg_4__2__10_ ( .D(n2961), .CK(clk), .RN(rst_n), .Q(
        w_matrix[474]) );
  DFFRHQX1 w_matrix_reg_4__6__10_ ( .D(n3025), .CK(clk), .RN(rst_n), .Q(
        w_matrix[410]) );
  DFFRHQX1 w_matrix_reg_5__2__10_ ( .D(n3089), .CK(clk), .RN(rst_n), .Q(
        w_matrix[346]) );
  DFFRHQX1 w_matrix_reg_5__6__10_ ( .D(n3153), .CK(clk), .RN(rst_n), .Q(
        w_matrix[282]) );
  DFFRHQX1 w_matrix_reg_6__2__10_ ( .D(n3217), .CK(clk), .RN(rst_n), .Q(
        w_matrix[218]) );
  DFFRHQX1 w_matrix_reg_6__6__10_ ( .D(n3281), .CK(clk), .RN(rst_n), .Q(
        w_matrix[154]) );
  DFFRHQX1 w_matrix_reg_7__2__10_ ( .D(n3345), .CK(clk), .RN(rst_n), .Q(
        w_matrix[90]) );
  DFFRHQX1 w_matrix_reg_7__6__10_ ( .D(n3409), .CK(clk), .RN(rst_n), .Q(
        w_matrix[26]) );
  DFFRHQX1 w_matrix_reg_1__2__9_ ( .D(n2578), .CK(clk), .RN(rst_n), .Q(
        w_matrix[857]) );
  DFFRHQX1 w_matrix_reg_1__6__9_ ( .D(n2642), .CK(clk), .RN(rst_n), .Q(
        w_matrix[793]) );
  DFFRHQX1 w_matrix_reg_2__2__9_ ( .D(n2706), .CK(clk), .RN(rst_n), .Q(
        w_matrix[729]) );
  DFFRHQX1 w_matrix_reg_2__6__9_ ( .D(n2770), .CK(clk), .RN(rst_n), .Q(
        w_matrix[665]) );
  DFFRHQX1 w_matrix_reg_3__2__9_ ( .D(n2834), .CK(clk), .RN(rst_n), .Q(
        w_matrix[601]) );
  DFFRHQX1 w_matrix_reg_3__6__9_ ( .D(n2898), .CK(clk), .RN(rst_n), .Q(
        w_matrix[537]) );
  DFFRHQX1 w_matrix_reg_4__2__9_ ( .D(n2962), .CK(clk), .RN(rst_n), .Q(
        w_matrix[473]) );
  DFFRHQX1 w_matrix_reg_4__6__9_ ( .D(n3026), .CK(clk), .RN(rst_n), .Q(
        w_matrix[409]) );
  DFFRHQX1 w_matrix_reg_5__2__9_ ( .D(n3090), .CK(clk), .RN(rst_n), .Q(
        w_matrix[345]) );
  DFFRHQX1 w_matrix_reg_5__6__9_ ( .D(n3154), .CK(clk), .RN(rst_n), .Q(
        w_matrix[281]) );
  DFFRHQX1 w_matrix_reg_6__2__9_ ( .D(n3218), .CK(clk), .RN(rst_n), .Q(
        w_matrix[217]) );
  DFFRHQX1 w_matrix_reg_6__6__9_ ( .D(n3282), .CK(clk), .RN(rst_n), .Q(
        w_matrix[153]) );
  DFFRHQX1 w_matrix_reg_7__2__9_ ( .D(n3346), .CK(clk), .RN(rst_n), .Q(
        w_matrix[89]) );
  DFFRHQX1 w_matrix_reg_7__6__9_ ( .D(n3410), .CK(clk), .RN(rst_n), .Q(
        w_matrix[25]) );
  DFFRHQX1 w_matrix_reg_1__2__8_ ( .D(n2579), .CK(clk), .RN(rst_n), .Q(
        w_matrix[856]) );
  DFFRHQX1 w_matrix_reg_1__6__8_ ( .D(n2643), .CK(clk), .RN(rst_n), .Q(
        w_matrix[792]) );
  DFFRHQX1 w_matrix_reg_2__2__8_ ( .D(n2707), .CK(clk), .RN(rst_n), .Q(
        w_matrix[728]) );
  DFFRHQX1 w_matrix_reg_2__6__8_ ( .D(n2771), .CK(clk), .RN(rst_n), .Q(
        w_matrix[664]) );
  DFFRHQX1 w_matrix_reg_3__2__8_ ( .D(n2835), .CK(clk), .RN(rst_n), .Q(
        w_matrix[600]) );
  DFFRHQX1 w_matrix_reg_3__6__8_ ( .D(n2899), .CK(clk), .RN(rst_n), .Q(
        w_matrix[536]) );
  DFFRHQX1 w_matrix_reg_4__2__8_ ( .D(n2963), .CK(clk), .RN(rst_n), .Q(
        w_matrix[472]) );
  DFFRHQX1 w_matrix_reg_4__6__8_ ( .D(n3027), .CK(clk), .RN(rst_n), .Q(
        w_matrix[408]) );
  DFFRHQX1 w_matrix_reg_5__2__8_ ( .D(n3091), .CK(clk), .RN(rst_n), .Q(
        w_matrix[344]) );
  DFFRHQX1 w_matrix_reg_5__6__8_ ( .D(n3155), .CK(clk), .RN(rst_n), .Q(
        w_matrix[280]) );
  DFFRHQX1 w_matrix_reg_6__2__8_ ( .D(n3219), .CK(clk), .RN(rst_n), .Q(
        w_matrix[216]) );
  DFFRHQX1 w_matrix_reg_6__6__8_ ( .D(n3283), .CK(clk), .RN(rst_n), .Q(
        w_matrix[152]) );
  DFFRHQX1 w_matrix_reg_7__2__8_ ( .D(n3347), .CK(clk), .RN(rst_n), .Q(
        w_matrix[88]) );
  DFFRHQX1 w_matrix_reg_7__6__8_ ( .D(n3411), .CK(clk), .RN(rst_n), .Q(
        w_matrix[24]) );
  DFFRHQX1 w_matrix_reg_1__3__10_ ( .D(n2593), .CK(clk), .RN(rst_n), .Q(
        w_matrix[842]) );
  DFFRHQX1 w_matrix_reg_1__7__10_ ( .D(n2657), .CK(clk), .RN(rst_n), .Q(
        w_matrix[778]) );
  DFFRHQX1 w_matrix_reg_2__3__10_ ( .D(n2721), .CK(clk), .RN(rst_n), .Q(
        w_matrix[714]) );
  DFFRHQX1 w_matrix_reg_2__7__10_ ( .D(n2785), .CK(clk), .RN(rst_n), .Q(
        w_matrix[650]) );
  DFFRHQX1 w_matrix_reg_3__3__10_ ( .D(n2849), .CK(clk), .RN(rst_n), .Q(
        w_matrix[586]) );
  DFFRHQX1 w_matrix_reg_3__7__10_ ( .D(n2913), .CK(clk), .RN(rst_n), .Q(
        w_matrix[522]) );
  DFFRHQX1 w_matrix_reg_4__3__10_ ( .D(n2977), .CK(clk), .RN(rst_n), .Q(
        w_matrix[458]) );
  DFFRHQX1 w_matrix_reg_4__7__10_ ( .D(n3041), .CK(clk), .RN(rst_n), .Q(
        w_matrix[394]) );
  DFFRHQX1 w_matrix_reg_5__3__10_ ( .D(n3105), .CK(clk), .RN(rst_n), .Q(
        w_matrix[330]) );
  DFFRHQX1 w_matrix_reg_5__7__10_ ( .D(n3169), .CK(clk), .RN(rst_n), .Q(
        w_matrix[266]) );
  DFFRHQX1 w_matrix_reg_6__3__10_ ( .D(n3233), .CK(clk), .RN(rst_n), .Q(
        w_matrix[202]) );
  DFFRHQX1 w_matrix_reg_6__7__10_ ( .D(n3297), .CK(clk), .RN(rst_n), .Q(
        w_matrix[138]) );
  DFFRHQX1 w_matrix_reg_7__3__10_ ( .D(n3361), .CK(clk), .RN(rst_n), .Q(
        w_matrix[74]) );
  DFFRHQX1 w_matrix_reg_7__7__10_ ( .D(n3425), .CK(clk), .RN(rst_n), .Q(
        w_matrix[10]) );
  DFFRX1 w_matrix_reg_1__1__7_ ( .D(n2564), .CK(clk), .RN(rst_n), .Q(
        w_matrix[871]), .QN(n666) );
  DFFRX1 w_matrix_reg_1__1__6_ ( .D(n2565), .CK(clk), .RN(rst_n), .Q(
        w_matrix[870]), .QN(n667) );
  DFFRX1 w_matrix_reg_1__1__5_ ( .D(n2566), .CK(clk), .RN(rst_n), .Q(
        w_matrix[869]), .QN(n668) );
  DFFRX1 w_matrix_reg_1__1__4_ ( .D(n2567), .CK(clk), .RN(rst_n), .Q(
        w_matrix[868]), .QN(n669) );
  DFFRX1 w_matrix_reg_1__1__3_ ( .D(n2568), .CK(clk), .RN(rst_n), .Q(
        w_matrix[867]), .QN(n670) );
  DFFRX1 w_matrix_reg_1__1__2_ ( .D(n2569), .CK(clk), .RN(rst_n), .Q(
        w_matrix[866]), .QN(n671) );
  DFFRX1 w_matrix_reg_1__1__1_ ( .D(n2570), .CK(clk), .RN(rst_n), .Q(
        w_matrix[865]), .QN(n672) );
  DFFRHQX1 inA41_reg_6_ ( .D(N11687), .CK(clk), .RN(rst_n), .Q(inA41[6]) );
  DFFRHQX1 inA81_reg_6_ ( .D(N12066), .CK(clk), .RN(rst_n), .Q(inA81[6]) );
  DFFRHQX1 inA51_reg_6_ ( .D(N11779), .CK(clk), .RN(rst_n), .Q(inA51[6]) );
  DFFRHQX1 inA51_reg_4_ ( .D(N11777), .CK(clk), .RN(rst_n), .Q(inA51[4]) );
  DFFRHQX1 inA51_reg_2_ ( .D(N11775), .CK(clk), .RN(rst_n), .Q(inA51[2]) );
  DFFRHQX1 inA41_reg_4_ ( .D(N11685), .CK(clk), .RN(rst_n), .Q(inA41[4]) );
  DFFRHQX1 inA81_reg_4_ ( .D(N12064), .CK(clk), .RN(rst_n), .Q(inA81[4]) );
  DFFRHQX1 inA21_reg_6_ ( .D(N11496), .CK(clk), .RN(rst_n), .Q(inA21[6]) );
  DFFRHQX1 inA61_reg_6_ ( .D(N11876), .CK(clk), .RN(rst_n), .Q(inA61[6]) );
  DFFRHQX1 inA21_reg_4_ ( .D(N11494), .CK(clk), .RN(rst_n), .Q(inA21[4]) );
  DFFRHQX1 inA61_reg_4_ ( .D(N11874), .CK(clk), .RN(rst_n), .Q(inA61[4]) );
  DFFRHQX1 inA61_reg_2_ ( .D(N11872), .CK(clk), .RN(rst_n), .Q(inA61[2]) );
  DFFRHQX1 inA21_reg_2_ ( .D(N11492), .CK(clk), .RN(rst_n), .Q(inA21[2]) );
  DFFRHQX1 inA41_reg_2_ ( .D(N11683), .CK(clk), .RN(rst_n), .Q(inA41[2]) );
  DFFRHQX1 inA81_reg_2_ ( .D(N12062), .CK(clk), .RN(rst_n), .Q(inA81[2]) );
  DFFRHQX1 inA31_reg_6_ ( .D(N11590), .CK(clk), .RN(rst_n), .Q(inA31[6]) );
  DFFRHQX1 inA71_reg_6_ ( .D(N11970), .CK(clk), .RN(rst_n), .Q(inA71[6]) );
  DFFRHQX1 inA31_reg_4_ ( .D(N11588), .CK(clk), .RN(rst_n), .Q(inA31[4]) );
  DFFRHQX1 inA71_reg_4_ ( .D(N11968), .CK(clk), .RN(rst_n), .Q(inA71[4]) );
  DFFRHQX1 inA31_reg_2_ ( .D(N11586), .CK(clk), .RN(rst_n), .Q(inA31[2]) );
  DFFRHQX1 inA71_reg_2_ ( .D(N11966), .CK(clk), .RN(rst_n), .Q(inA71[2]) );
  DFFRHQX1 inA41_reg_7_ ( .D(N11688), .CK(clk), .RN(rst_n), .Q(inA41[7]) );
  DFFRHQX1 inA81_reg_7_ ( .D(N12067), .CK(clk), .RN(rst_n), .Q(inA81[7]) );
  DFFRHQX1 inA41_reg_5_ ( .D(N11686), .CK(clk), .RN(rst_n), .Q(inA41[5]) );
  DFFRHQX1 inA81_reg_5_ ( .D(N12065), .CK(clk), .RN(rst_n), .Q(inA81[5]) );
  DFFRHQX1 inA51_reg_7_ ( .D(N11780), .CK(clk), .RN(rst_n), .Q(inA51[7]) );
  DFFRHQX1 inA51_reg_5_ ( .D(N11778), .CK(clk), .RN(rst_n), .Q(inA51[5]) );
  DFFRHQX1 inA51_reg_3_ ( .D(N11776), .CK(clk), .RN(rst_n), .Q(inA51[3]) );
  DFFRHQX1 inA41_reg_3_ ( .D(N11684), .CK(clk), .RN(rst_n), .Q(inA41[3]) );
  DFFRHQX1 inA81_reg_3_ ( .D(N12063), .CK(clk), .RN(rst_n), .Q(inA81[3]) );
  DFFRHQX1 inA21_reg_7_ ( .D(N11497), .CK(clk), .RN(rst_n), .Q(inA21[7]) );
  DFFRHQX1 inA61_reg_7_ ( .D(N11877), .CK(clk), .RN(rst_n), .Q(inA61[7]) );
  DFFRHQX1 inA21_reg_5_ ( .D(N11495), .CK(clk), .RN(rst_n), .Q(inA21[5]) );
  DFFRHQX1 inA61_reg_5_ ( .D(N11875), .CK(clk), .RN(rst_n), .Q(inA61[5]) );
  DFFRHQX1 inA21_reg_3_ ( .D(N11493), .CK(clk), .RN(rst_n), .Q(inA21[3]) );
  DFFRHQX1 inA61_reg_3_ ( .D(N11873), .CK(clk), .RN(rst_n), .Q(inA61[3]) );
  DFFRHQX1 inA31_reg_7_ ( .D(N11591), .CK(clk), .RN(rst_n), .Q(inA31[7]) );
  DFFRHQX1 inA71_reg_7_ ( .D(N11971), .CK(clk), .RN(rst_n), .Q(inA71[7]) );
  DFFRHQX1 inA31_reg_5_ ( .D(N11589), .CK(clk), .RN(rst_n), .Q(inA31[5]) );
  DFFRHQX1 inA71_reg_5_ ( .D(N11969), .CK(clk), .RN(rst_n), .Q(inA71[5]) );
  DFFRHQX1 inA31_reg_3_ ( .D(N11587), .CK(clk), .RN(rst_n), .Q(inA31[3]) );
  DFFRHQX1 inA71_reg_3_ ( .D(N11967), .CK(clk), .RN(rst_n), .Q(inA71[3]) );
  DFFRHQX1 w_matrix_reg_1__4__0_ ( .D(n2619), .CK(clk), .RN(rst_n), .Q(
        w_matrix[816]) );
  DFFRHQX1 w_matrix_reg_2__0__0_ ( .D(n2683), .CK(clk), .RN(rst_n), .Q(
        w_matrix[752]) );
  DFFRHQX1 w_matrix_reg_2__4__0_ ( .D(n2747), .CK(clk), .RN(rst_n), .Q(
        w_matrix[688]) );
  DFFRHQX1 w_matrix_reg_3__0__0_ ( .D(n2811), .CK(clk), .RN(rst_n), .Q(
        w_matrix[624]) );
  DFFRHQX1 w_matrix_reg_3__4__0_ ( .D(n2875), .CK(clk), .RN(rst_n), .Q(
        w_matrix[560]) );
  DFFRHQX1 w_matrix_reg_4__0__0_ ( .D(n2939), .CK(clk), .RN(rst_n), .Q(
        w_matrix[496]) );
  DFFRHQX1 w_matrix_reg_4__4__0_ ( .D(n3003), .CK(clk), .RN(rst_n), .Q(
        w_matrix[432]) );
  DFFRHQX1 w_matrix_reg_5__0__0_ ( .D(n3067), .CK(clk), .RN(rst_n), .Q(
        w_matrix[368]) );
  DFFRHQX1 w_matrix_reg_5__4__0_ ( .D(n3131), .CK(clk), .RN(rst_n), .Q(
        w_matrix[304]) );
  DFFRHQX1 w_matrix_reg_6__0__0_ ( .D(n3195), .CK(clk), .RN(rst_n), .Q(
        w_matrix[240]) );
  DFFRHQX1 w_matrix_reg_6__4__0_ ( .D(n3259), .CK(clk), .RN(rst_n), .Q(
        w_matrix[176]) );
  DFFRHQX1 w_matrix_reg_7__0__0_ ( .D(n3323), .CK(clk), .RN(rst_n), .Q(
        w_matrix[112]) );
  DFFRHQX1 w_matrix_reg_7__4__0_ ( .D(n3387), .CK(clk), .RN(rst_n), .Q(
        w_matrix[48]) );
  DFFRHQX1 w_matrix_reg_1__5__0_ ( .D(n2635), .CK(clk), .RN(rst_n), .Q(
        w_matrix[800]) );
  DFFRHQX1 w_matrix_reg_2__1__0_ ( .D(n2699), .CK(clk), .RN(rst_n), .Q(
        w_matrix[736]) );
  DFFRHQX1 w_matrix_reg_2__5__0_ ( .D(n2763), .CK(clk), .RN(rst_n), .Q(
        w_matrix[672]) );
  DFFRHQX1 w_matrix_reg_3__1__0_ ( .D(n2827), .CK(clk), .RN(rst_n), .Q(
        w_matrix[608]) );
  DFFRHQX1 w_matrix_reg_3__5__0_ ( .D(n2891), .CK(clk), .RN(rst_n), .Q(
        w_matrix[544]) );
  DFFRHQX1 w_matrix_reg_4__1__0_ ( .D(n2955), .CK(clk), .RN(rst_n), .Q(
        w_matrix[480]) );
  DFFRHQX1 w_matrix_reg_4__5__0_ ( .D(n3019), .CK(clk), .RN(rst_n), .Q(
        w_matrix[416]) );
  DFFRHQX1 w_matrix_reg_5__1__0_ ( .D(n3083), .CK(clk), .RN(rst_n), .Q(
        w_matrix[352]) );
  DFFRHQX1 w_matrix_reg_5__5__0_ ( .D(n3147), .CK(clk), .RN(rst_n), .Q(
        w_matrix[288]) );
  DFFRHQX1 w_matrix_reg_6__1__0_ ( .D(n3211), .CK(clk), .RN(rst_n), .Q(
        w_matrix[224]) );
  DFFRHQX1 w_matrix_reg_6__5__0_ ( .D(n3275), .CK(clk), .RN(rst_n), .Q(
        w_matrix[160]) );
  DFFRHQX1 w_matrix_reg_7__1__0_ ( .D(n3339), .CK(clk), .RN(rst_n), .Q(
        w_matrix[96]) );
  DFFRHQX1 w_matrix_reg_7__5__0_ ( .D(n3403), .CK(clk), .RN(rst_n), .Q(
        w_matrix[32]) );
  DFFRHQX1 w_matrix_reg_1__2__0_ ( .D(n2587), .CK(clk), .RN(rst_n), .Q(
        w_matrix[848]) );
  DFFRHQX1 w_matrix_reg_1__6__0_ ( .D(n2651), .CK(clk), .RN(rst_n), .Q(
        w_matrix[784]) );
  DFFRHQX1 w_matrix_reg_2__2__0_ ( .D(n2715), .CK(clk), .RN(rst_n), .Q(
        w_matrix[720]) );
  DFFRHQX1 w_matrix_reg_2__6__0_ ( .D(n2779), .CK(clk), .RN(rst_n), .Q(
        w_matrix[656]) );
  DFFRHQX1 w_matrix_reg_3__2__0_ ( .D(n2843), .CK(clk), .RN(rst_n), .Q(
        w_matrix[592]) );
  DFFRHQX1 w_matrix_reg_3__6__0_ ( .D(n2907), .CK(clk), .RN(rst_n), .Q(
        w_matrix[528]) );
  DFFRHQX1 w_matrix_reg_4__2__0_ ( .D(n2971), .CK(clk), .RN(rst_n), .Q(
        w_matrix[464]) );
  DFFRHQX1 w_matrix_reg_4__6__0_ ( .D(n3035), .CK(clk), .RN(rst_n), .Q(
        w_matrix[400]) );
  DFFRHQX1 w_matrix_reg_5__2__0_ ( .D(n3099), .CK(clk), .RN(rst_n), .Q(
        w_matrix[336]) );
  DFFRHQX1 w_matrix_reg_5__6__0_ ( .D(n3163), .CK(clk), .RN(rst_n), .Q(
        w_matrix[272]) );
  DFFRHQX1 w_matrix_reg_6__2__0_ ( .D(n3227), .CK(clk), .RN(rst_n), .Q(
        w_matrix[208]) );
  DFFRHQX1 w_matrix_reg_6__6__0_ ( .D(n3291), .CK(clk), .RN(rst_n), .Q(
        w_matrix[144]) );
  DFFRHQX1 w_matrix_reg_7__2__0_ ( .D(n3355), .CK(clk), .RN(rst_n), .Q(
        w_matrix[80]) );
  DFFRHQX1 w_matrix_reg_7__6__0_ ( .D(n3419), .CK(clk), .RN(rst_n), .Q(
        w_matrix[16]) );
  DFFRHQX1 w_matrix_reg_1__3__0_ ( .D(n2603), .CK(clk), .RN(rst_n), .Q(
        w_matrix[832]) );
  DFFRHQX1 w_matrix_reg_1__7__0_ ( .D(n2667), .CK(clk), .RN(rst_n), .Q(
        w_matrix[768]) );
  DFFRHQX1 w_matrix_reg_2__3__0_ ( .D(n2731), .CK(clk), .RN(rst_n), .Q(
        w_matrix[704]) );
  DFFRHQX1 w_matrix_reg_2__7__0_ ( .D(n2795), .CK(clk), .RN(rst_n), .Q(
        w_matrix[640]) );
  DFFRHQX1 w_matrix_reg_3__3__0_ ( .D(n2859), .CK(clk), .RN(rst_n), .Q(
        w_matrix[576]) );
  DFFRHQX1 w_matrix_reg_3__7__0_ ( .D(n2923), .CK(clk), .RN(rst_n), .Q(
        w_matrix[512]) );
  DFFRHQX1 w_matrix_reg_4__3__0_ ( .D(n2987), .CK(clk), .RN(rst_n), .Q(
        w_matrix[448]) );
  DFFRHQX1 w_matrix_reg_4__7__0_ ( .D(n3051), .CK(clk), .RN(rst_n), .Q(
        w_matrix[384]) );
  DFFRHQX1 w_matrix_reg_5__3__0_ ( .D(n3115), .CK(clk), .RN(rst_n), .Q(
        w_matrix[320]) );
  DFFRHQX1 w_matrix_reg_5__7__0_ ( .D(n3179), .CK(clk), .RN(rst_n), .Q(
        w_matrix[256]) );
  DFFRHQX1 w_matrix_reg_6__3__0_ ( .D(n3243), .CK(clk), .RN(rst_n), .Q(
        w_matrix[192]) );
  DFFRHQX1 w_matrix_reg_6__7__0_ ( .D(n3307), .CK(clk), .RN(rst_n), .Q(
        w_matrix[128]) );
  DFFRHQX1 w_matrix_reg_7__3__0_ ( .D(n3371), .CK(clk), .RN(rst_n), .Q(
        w_matrix[64]) );
  DFFRHQX1 w_matrix_reg_7__7__0_ ( .D(n3435), .CK(clk), .RN(rst_n), .Q(
        w_matrix[0]) );
  DFFRHQX1 w_matrix_reg_1__3__7_ ( .D(n2596), .CK(clk), .RN(rst_n), .Q(
        w_matrix[839]) );
  DFFRHQX1 w_matrix_reg_1__7__7_ ( .D(n2660), .CK(clk), .RN(rst_n), .Q(
        w_matrix[775]) );
  DFFRHQX1 w_matrix_reg_2__3__7_ ( .D(n2724), .CK(clk), .RN(rst_n), .Q(
        w_matrix[711]) );
  DFFRHQX1 w_matrix_reg_2__7__7_ ( .D(n2788), .CK(clk), .RN(rst_n), .Q(
        w_matrix[647]) );
  DFFRHQX1 w_matrix_reg_3__3__7_ ( .D(n2852), .CK(clk), .RN(rst_n), .Q(
        w_matrix[583]) );
  DFFRHQX1 w_matrix_reg_3__7__7_ ( .D(n2916), .CK(clk), .RN(rst_n), .Q(
        w_matrix[519]) );
  DFFRHQX1 w_matrix_reg_4__3__7_ ( .D(n2980), .CK(clk), .RN(rst_n), .Q(
        w_matrix[455]) );
  DFFRHQX1 w_matrix_reg_4__7__7_ ( .D(n3044), .CK(clk), .RN(rst_n), .Q(
        w_matrix[391]) );
  DFFRHQX1 w_matrix_reg_5__3__7_ ( .D(n3108), .CK(clk), .RN(rst_n), .Q(
        w_matrix[327]) );
  DFFRHQX1 w_matrix_reg_5__7__7_ ( .D(n3172), .CK(clk), .RN(rst_n), .Q(
        w_matrix[263]) );
  DFFRHQX1 w_matrix_reg_6__3__7_ ( .D(n3236), .CK(clk), .RN(rst_n), .Q(
        w_matrix[199]) );
  DFFRHQX1 w_matrix_reg_6__7__7_ ( .D(n3300), .CK(clk), .RN(rst_n), .Q(
        w_matrix[135]) );
  DFFRHQX1 w_matrix_reg_7__3__7_ ( .D(n3364), .CK(clk), .RN(rst_n), .Q(
        w_matrix[71]) );
  DFFRHQX1 w_matrix_reg_7__7__7_ ( .D(n3428), .CK(clk), .RN(rst_n), .Q(
        w_matrix[7]) );
  DFFRHQX1 w_matrix_reg_1__3__6_ ( .D(n2597), .CK(clk), .RN(rst_n), .Q(
        w_matrix[838]) );
  DFFRHQX1 w_matrix_reg_1__7__6_ ( .D(n2661), .CK(clk), .RN(rst_n), .Q(
        w_matrix[774]) );
  DFFRHQX1 w_matrix_reg_2__3__6_ ( .D(n2725), .CK(clk), .RN(rst_n), .Q(
        w_matrix[710]) );
  DFFRHQX1 w_matrix_reg_2__7__6_ ( .D(n2789), .CK(clk), .RN(rst_n), .Q(
        w_matrix[646]) );
  DFFRHQX1 w_matrix_reg_3__3__6_ ( .D(n2853), .CK(clk), .RN(rst_n), .Q(
        w_matrix[582]) );
  DFFRHQX1 w_matrix_reg_3__7__6_ ( .D(n2917), .CK(clk), .RN(rst_n), .Q(
        w_matrix[518]) );
  DFFRHQX1 w_matrix_reg_4__3__6_ ( .D(n2981), .CK(clk), .RN(rst_n), .Q(
        w_matrix[454]) );
  DFFRHQX1 w_matrix_reg_4__7__6_ ( .D(n3045), .CK(clk), .RN(rst_n), .Q(
        w_matrix[390]) );
  DFFRHQX1 w_matrix_reg_5__3__6_ ( .D(n3109), .CK(clk), .RN(rst_n), .Q(
        w_matrix[326]) );
  DFFRHQX1 w_matrix_reg_5__7__6_ ( .D(n3173), .CK(clk), .RN(rst_n), .Q(
        w_matrix[262]) );
  DFFRHQX1 w_matrix_reg_6__3__6_ ( .D(n3237), .CK(clk), .RN(rst_n), .Q(
        w_matrix[198]) );
  DFFRHQX1 w_matrix_reg_6__7__6_ ( .D(n3301), .CK(clk), .RN(rst_n), .Q(
        w_matrix[134]) );
  DFFRHQX1 w_matrix_reg_7__3__6_ ( .D(n3365), .CK(clk), .RN(rst_n), .Q(
        w_matrix[70]) );
  DFFRHQX1 w_matrix_reg_7__7__6_ ( .D(n3429), .CK(clk), .RN(rst_n), .Q(
        w_matrix[6]) );
  DFFRHQX1 w_matrix_reg_1__3__5_ ( .D(n2598), .CK(clk), .RN(rst_n), .Q(
        w_matrix[837]) );
  DFFRHQX1 w_matrix_reg_1__7__5_ ( .D(n2662), .CK(clk), .RN(rst_n), .Q(
        w_matrix[773]) );
  DFFRHQX1 w_matrix_reg_2__3__5_ ( .D(n2726), .CK(clk), .RN(rst_n), .Q(
        w_matrix[709]) );
  DFFRHQX1 w_matrix_reg_2__7__5_ ( .D(n2790), .CK(clk), .RN(rst_n), .Q(
        w_matrix[645]) );
  DFFRHQX1 w_matrix_reg_3__3__5_ ( .D(n2854), .CK(clk), .RN(rst_n), .Q(
        w_matrix[581]) );
  DFFRHQX1 w_matrix_reg_3__7__5_ ( .D(n2918), .CK(clk), .RN(rst_n), .Q(
        w_matrix[517]) );
  DFFRHQX1 w_matrix_reg_4__3__5_ ( .D(n2982), .CK(clk), .RN(rst_n), .Q(
        w_matrix[453]) );
  DFFRHQX1 w_matrix_reg_4__7__5_ ( .D(n3046), .CK(clk), .RN(rst_n), .Q(
        w_matrix[389]) );
  DFFRHQX1 w_matrix_reg_5__3__5_ ( .D(n3110), .CK(clk), .RN(rst_n), .Q(
        w_matrix[325]) );
  DFFRHQX1 w_matrix_reg_5__7__5_ ( .D(n3174), .CK(clk), .RN(rst_n), .Q(
        w_matrix[261]) );
  DFFRHQX1 w_matrix_reg_6__3__5_ ( .D(n3238), .CK(clk), .RN(rst_n), .Q(
        w_matrix[197]) );
  DFFRHQX1 w_matrix_reg_6__7__5_ ( .D(n3302), .CK(clk), .RN(rst_n), .Q(
        w_matrix[133]) );
  DFFRHQX1 w_matrix_reg_7__3__5_ ( .D(n3366), .CK(clk), .RN(rst_n), .Q(
        w_matrix[69]) );
  DFFRHQX1 w_matrix_reg_7__7__5_ ( .D(n3430), .CK(clk), .RN(rst_n), .Q(
        w_matrix[5]) );
  DFFRHQX1 w_matrix_reg_1__4__7_ ( .D(n2612), .CK(clk), .RN(rst_n), .Q(
        w_matrix[823]) );
  DFFRHQX1 w_matrix_reg_2__0__7_ ( .D(n2676), .CK(clk), .RN(rst_n), .Q(
        w_matrix[759]) );
  DFFRHQX1 w_matrix_reg_2__4__7_ ( .D(n2740), .CK(clk), .RN(rst_n), .Q(
        w_matrix[695]) );
  DFFRHQX1 w_matrix_reg_3__0__7_ ( .D(n2804), .CK(clk), .RN(rst_n), .Q(
        w_matrix[631]) );
  DFFRHQX1 w_matrix_reg_3__4__7_ ( .D(n2868), .CK(clk), .RN(rst_n), .Q(
        w_matrix[567]) );
  DFFRHQX1 w_matrix_reg_4__0__7_ ( .D(n2932), .CK(clk), .RN(rst_n), .Q(
        w_matrix[503]) );
  DFFRHQX1 w_matrix_reg_4__4__7_ ( .D(n2996), .CK(clk), .RN(rst_n), .Q(
        w_matrix[439]) );
  DFFRHQX1 w_matrix_reg_5__0__7_ ( .D(n3060), .CK(clk), .RN(rst_n), .Q(
        w_matrix[375]) );
  DFFRHQX1 w_matrix_reg_5__4__7_ ( .D(n3124), .CK(clk), .RN(rst_n), .Q(
        w_matrix[311]) );
  DFFRHQX1 w_matrix_reg_6__0__7_ ( .D(n3188), .CK(clk), .RN(rst_n), .Q(
        w_matrix[247]) );
  DFFRHQX1 w_matrix_reg_6__4__7_ ( .D(n3252), .CK(clk), .RN(rst_n), .Q(
        w_matrix[183]) );
  DFFRHQX1 w_matrix_reg_7__0__7_ ( .D(n3316), .CK(clk), .RN(rst_n), .Q(
        w_matrix[119]) );
  DFFRHQX1 w_matrix_reg_7__4__7_ ( .D(n3380), .CK(clk), .RN(rst_n), .Q(
        w_matrix[55]) );
  DFFRHQX1 w_matrix_reg_1__4__6_ ( .D(n2613), .CK(clk), .RN(rst_n), .Q(
        w_matrix[822]) );
  DFFRHQX1 w_matrix_reg_2__0__6_ ( .D(n2677), .CK(clk), .RN(rst_n), .Q(
        w_matrix[758]) );
  DFFRHQX1 w_matrix_reg_2__4__6_ ( .D(n2741), .CK(clk), .RN(rst_n), .Q(
        w_matrix[694]) );
  DFFRHQX1 w_matrix_reg_3__0__6_ ( .D(n2805), .CK(clk), .RN(rst_n), .Q(
        w_matrix[630]) );
  DFFRHQX1 w_matrix_reg_3__4__6_ ( .D(n2869), .CK(clk), .RN(rst_n), .Q(
        w_matrix[566]) );
  DFFRHQX1 w_matrix_reg_4__0__6_ ( .D(n2933), .CK(clk), .RN(rst_n), .Q(
        w_matrix[502]) );
  DFFRHQX1 w_matrix_reg_4__4__6_ ( .D(n2997), .CK(clk), .RN(rst_n), .Q(
        w_matrix[438]) );
  DFFRHQX1 w_matrix_reg_5__0__6_ ( .D(n3061), .CK(clk), .RN(rst_n), .Q(
        w_matrix[374]) );
  DFFRHQX1 w_matrix_reg_5__4__6_ ( .D(n3125), .CK(clk), .RN(rst_n), .Q(
        w_matrix[310]) );
  DFFRHQX1 w_matrix_reg_6__0__6_ ( .D(n3189), .CK(clk), .RN(rst_n), .Q(
        w_matrix[246]) );
  DFFRHQX1 w_matrix_reg_6__4__6_ ( .D(n3253), .CK(clk), .RN(rst_n), .Q(
        w_matrix[182]) );
  DFFRHQX1 w_matrix_reg_7__0__6_ ( .D(n3317), .CK(clk), .RN(rst_n), .Q(
        w_matrix[118]) );
  DFFRHQX1 w_matrix_reg_7__4__6_ ( .D(n3381), .CK(clk), .RN(rst_n), .Q(
        w_matrix[54]) );
  DFFRHQX1 w_matrix_reg_1__4__5_ ( .D(n2614), .CK(clk), .RN(rst_n), .Q(
        w_matrix[821]) );
  DFFRHQX1 w_matrix_reg_2__0__5_ ( .D(n2678), .CK(clk), .RN(rst_n), .Q(
        w_matrix[757]) );
  DFFRHQX1 w_matrix_reg_2__4__5_ ( .D(n2742), .CK(clk), .RN(rst_n), .Q(
        w_matrix[693]) );
  DFFRHQX1 w_matrix_reg_3__0__5_ ( .D(n2806), .CK(clk), .RN(rst_n), .Q(
        w_matrix[629]) );
  DFFRHQX1 w_matrix_reg_3__4__5_ ( .D(n2870), .CK(clk), .RN(rst_n), .Q(
        w_matrix[565]) );
  DFFRHQX1 w_matrix_reg_4__0__5_ ( .D(n2934), .CK(clk), .RN(rst_n), .Q(
        w_matrix[501]) );
  DFFRHQX1 w_matrix_reg_4__4__5_ ( .D(n2998), .CK(clk), .RN(rst_n), .Q(
        w_matrix[437]) );
  DFFRHQX1 w_matrix_reg_5__0__5_ ( .D(n3062), .CK(clk), .RN(rst_n), .Q(
        w_matrix[373]) );
  DFFRHQX1 w_matrix_reg_5__4__5_ ( .D(n3126), .CK(clk), .RN(rst_n), .Q(
        w_matrix[309]) );
  DFFRHQX1 w_matrix_reg_6__0__5_ ( .D(n3190), .CK(clk), .RN(rst_n), .Q(
        w_matrix[245]) );
  DFFRHQX1 w_matrix_reg_6__4__5_ ( .D(n3254), .CK(clk), .RN(rst_n), .Q(
        w_matrix[181]) );
  DFFRHQX1 w_matrix_reg_7__0__5_ ( .D(n3318), .CK(clk), .RN(rst_n), .Q(
        w_matrix[117]) );
  DFFRHQX1 w_matrix_reg_7__4__5_ ( .D(n3382), .CK(clk), .RN(rst_n), .Q(
        w_matrix[53]) );
  DFFRHQX1 w_matrix_reg_1__4__4_ ( .D(n2615), .CK(clk), .RN(rst_n), .Q(
        w_matrix[820]) );
  DFFRHQX1 w_matrix_reg_2__0__4_ ( .D(n2679), .CK(clk), .RN(rst_n), .Q(
        w_matrix[756]) );
  DFFRHQX1 w_matrix_reg_2__4__4_ ( .D(n2743), .CK(clk), .RN(rst_n), .Q(
        w_matrix[692]) );
  DFFRHQX1 w_matrix_reg_3__0__4_ ( .D(n2807), .CK(clk), .RN(rst_n), .Q(
        w_matrix[628]) );
  DFFRHQX1 w_matrix_reg_3__4__4_ ( .D(n2871), .CK(clk), .RN(rst_n), .Q(
        w_matrix[564]) );
  DFFRHQX1 w_matrix_reg_4__0__4_ ( .D(n2935), .CK(clk), .RN(rst_n), .Q(
        w_matrix[500]) );
  DFFRHQX1 w_matrix_reg_4__4__4_ ( .D(n2999), .CK(clk), .RN(rst_n), .Q(
        w_matrix[436]) );
  DFFRHQX1 w_matrix_reg_5__0__4_ ( .D(n3063), .CK(clk), .RN(rst_n), .Q(
        w_matrix[372]) );
  DFFRHQX1 w_matrix_reg_5__4__4_ ( .D(n3127), .CK(clk), .RN(rst_n), .Q(
        w_matrix[308]) );
  DFFRHQX1 w_matrix_reg_6__0__4_ ( .D(n3191), .CK(clk), .RN(rst_n), .Q(
        w_matrix[244]) );
  DFFRHQX1 w_matrix_reg_6__4__4_ ( .D(n3255), .CK(clk), .RN(rst_n), .Q(
        w_matrix[180]) );
  DFFRHQX1 w_matrix_reg_7__0__4_ ( .D(n3319), .CK(clk), .RN(rst_n), .Q(
        w_matrix[116]) );
  DFFRHQX1 w_matrix_reg_7__4__4_ ( .D(n3383), .CK(clk), .RN(rst_n), .Q(
        w_matrix[52]) );
  DFFRHQX1 w_matrix_reg_1__4__3_ ( .D(n2616), .CK(clk), .RN(rst_n), .Q(
        w_matrix[819]) );
  DFFRHQX1 w_matrix_reg_2__0__3_ ( .D(n2680), .CK(clk), .RN(rst_n), .Q(
        w_matrix[755]) );
  DFFRHQX1 w_matrix_reg_2__4__3_ ( .D(n2744), .CK(clk), .RN(rst_n), .Q(
        w_matrix[691]) );
  DFFRHQX1 w_matrix_reg_3__0__3_ ( .D(n2808), .CK(clk), .RN(rst_n), .Q(
        w_matrix[627]) );
  DFFRHQX1 w_matrix_reg_3__4__3_ ( .D(n2872), .CK(clk), .RN(rst_n), .Q(
        w_matrix[563]) );
  DFFRHQX1 w_matrix_reg_4__0__3_ ( .D(n2936), .CK(clk), .RN(rst_n), .Q(
        w_matrix[499]) );
  DFFRHQX1 w_matrix_reg_4__4__3_ ( .D(n3000), .CK(clk), .RN(rst_n), .Q(
        w_matrix[435]) );
  DFFRHQX1 w_matrix_reg_5__0__3_ ( .D(n3064), .CK(clk), .RN(rst_n), .Q(
        w_matrix[371]) );
  DFFRHQX1 w_matrix_reg_5__4__3_ ( .D(n3128), .CK(clk), .RN(rst_n), .Q(
        w_matrix[307]) );
  DFFRHQX1 w_matrix_reg_6__0__3_ ( .D(n3192), .CK(clk), .RN(rst_n), .Q(
        w_matrix[243]) );
  DFFRHQX1 w_matrix_reg_6__4__3_ ( .D(n3256), .CK(clk), .RN(rst_n), .Q(
        w_matrix[179]) );
  DFFRHQX1 w_matrix_reg_7__0__3_ ( .D(n3320), .CK(clk), .RN(rst_n), .Q(
        w_matrix[115]) );
  DFFRHQX1 w_matrix_reg_7__4__3_ ( .D(n3384), .CK(clk), .RN(rst_n), .Q(
        w_matrix[51]) );
  DFFRHQX1 w_matrix_reg_1__4__2_ ( .D(n2617), .CK(clk), .RN(rst_n), .Q(
        w_matrix[818]) );
  DFFRHQX1 w_matrix_reg_2__0__2_ ( .D(n2681), .CK(clk), .RN(rst_n), .Q(
        w_matrix[754]) );
  DFFRHQX1 w_matrix_reg_2__4__2_ ( .D(n2745), .CK(clk), .RN(rst_n), .Q(
        w_matrix[690]) );
  DFFRHQX1 w_matrix_reg_3__0__2_ ( .D(n2809), .CK(clk), .RN(rst_n), .Q(
        w_matrix[626]) );
  DFFRHQX1 w_matrix_reg_3__4__2_ ( .D(n2873), .CK(clk), .RN(rst_n), .Q(
        w_matrix[562]) );
  DFFRHQX1 w_matrix_reg_4__0__2_ ( .D(n2937), .CK(clk), .RN(rst_n), .Q(
        w_matrix[498]) );
  DFFRHQX1 w_matrix_reg_4__4__2_ ( .D(n3001), .CK(clk), .RN(rst_n), .Q(
        w_matrix[434]) );
  DFFRHQX1 w_matrix_reg_5__0__2_ ( .D(n3065), .CK(clk), .RN(rst_n), .Q(
        w_matrix[370]) );
  DFFRHQX1 w_matrix_reg_5__4__2_ ( .D(n3129), .CK(clk), .RN(rst_n), .Q(
        w_matrix[306]) );
  DFFRHQX1 w_matrix_reg_6__0__2_ ( .D(n3193), .CK(clk), .RN(rst_n), .Q(
        w_matrix[242]) );
  DFFRHQX1 w_matrix_reg_6__4__2_ ( .D(n3257), .CK(clk), .RN(rst_n), .Q(
        w_matrix[178]) );
  DFFRHQX1 w_matrix_reg_7__0__2_ ( .D(n3321), .CK(clk), .RN(rst_n), .Q(
        w_matrix[114]) );
  DFFRHQX1 w_matrix_reg_7__4__2_ ( .D(n3385), .CK(clk), .RN(rst_n), .Q(
        w_matrix[50]) );
  DFFRHQX1 w_matrix_reg_1__3__4_ ( .D(n2599), .CK(clk), .RN(rst_n), .Q(
        w_matrix[836]) );
  DFFRHQX1 w_matrix_reg_1__7__4_ ( .D(n2663), .CK(clk), .RN(rst_n), .Q(
        w_matrix[772]) );
  DFFRHQX1 w_matrix_reg_2__3__4_ ( .D(n2727), .CK(clk), .RN(rst_n), .Q(
        w_matrix[708]) );
  DFFRHQX1 w_matrix_reg_2__7__4_ ( .D(n2791), .CK(clk), .RN(rst_n), .Q(
        w_matrix[644]) );
  DFFRHQX1 w_matrix_reg_3__3__4_ ( .D(n2855), .CK(clk), .RN(rst_n), .Q(
        w_matrix[580]) );
  DFFRHQX1 w_matrix_reg_3__7__4_ ( .D(n2919), .CK(clk), .RN(rst_n), .Q(
        w_matrix[516]) );
  DFFRHQX1 w_matrix_reg_4__3__4_ ( .D(n2983), .CK(clk), .RN(rst_n), .Q(
        w_matrix[452]) );
  DFFRHQX1 w_matrix_reg_4__7__4_ ( .D(n3047), .CK(clk), .RN(rst_n), .Q(
        w_matrix[388]) );
  DFFRHQX1 w_matrix_reg_5__3__4_ ( .D(n3111), .CK(clk), .RN(rst_n), .Q(
        w_matrix[324]) );
  DFFRHQX1 w_matrix_reg_5__7__4_ ( .D(n3175), .CK(clk), .RN(rst_n), .Q(
        w_matrix[260]) );
  DFFRHQX1 w_matrix_reg_6__3__4_ ( .D(n3239), .CK(clk), .RN(rst_n), .Q(
        w_matrix[196]) );
  DFFRHQX1 w_matrix_reg_6__7__4_ ( .D(n3303), .CK(clk), .RN(rst_n), .Q(
        w_matrix[132]) );
  DFFRHQX1 w_matrix_reg_7__3__4_ ( .D(n3367), .CK(clk), .RN(rst_n), .Q(
        w_matrix[68]) );
  DFFRHQX1 w_matrix_reg_7__7__4_ ( .D(n3431), .CK(clk), .RN(rst_n), .Q(
        w_matrix[4]) );
  DFFRHQX1 w_matrix_reg_1__4__1_ ( .D(n2618), .CK(clk), .RN(rst_n), .Q(
        w_matrix[817]) );
  DFFRHQX1 w_matrix_reg_2__0__1_ ( .D(n2682), .CK(clk), .RN(rst_n), .Q(
        w_matrix[753]) );
  DFFRHQX1 w_matrix_reg_2__4__1_ ( .D(n2746), .CK(clk), .RN(rst_n), .Q(
        w_matrix[689]) );
  DFFRHQX1 w_matrix_reg_3__0__1_ ( .D(n2810), .CK(clk), .RN(rst_n), .Q(
        w_matrix[625]) );
  DFFRHQX1 w_matrix_reg_3__4__1_ ( .D(n2874), .CK(clk), .RN(rst_n), .Q(
        w_matrix[561]) );
  DFFRHQX1 w_matrix_reg_4__0__1_ ( .D(n2938), .CK(clk), .RN(rst_n), .Q(
        w_matrix[497]) );
  DFFRHQX1 w_matrix_reg_4__4__1_ ( .D(n3002), .CK(clk), .RN(rst_n), .Q(
        w_matrix[433]) );
  DFFRHQX1 w_matrix_reg_5__0__1_ ( .D(n3066), .CK(clk), .RN(rst_n), .Q(
        w_matrix[369]) );
  DFFRHQX1 w_matrix_reg_5__4__1_ ( .D(n3130), .CK(clk), .RN(rst_n), .Q(
        w_matrix[305]) );
  DFFRHQX1 w_matrix_reg_6__0__1_ ( .D(n3194), .CK(clk), .RN(rst_n), .Q(
        w_matrix[241]) );
  DFFRHQX1 w_matrix_reg_6__4__1_ ( .D(n3258), .CK(clk), .RN(rst_n), .Q(
        w_matrix[177]) );
  DFFRHQX1 w_matrix_reg_7__0__1_ ( .D(n3322), .CK(clk), .RN(rst_n), .Q(
        w_matrix[113]) );
  DFFRHQX1 w_matrix_reg_7__4__1_ ( .D(n3386), .CK(clk), .RN(rst_n), .Q(
        w_matrix[49]) );
  DFFRHQX1 w_matrix_reg_1__3__3_ ( .D(n2600), .CK(clk), .RN(rst_n), .Q(
        w_matrix[835]) );
  DFFRHQX1 w_matrix_reg_1__7__3_ ( .D(n2664), .CK(clk), .RN(rst_n), .Q(
        w_matrix[771]) );
  DFFRHQX1 w_matrix_reg_2__3__3_ ( .D(n2728), .CK(clk), .RN(rst_n), .Q(
        w_matrix[707]) );
  DFFRHQX1 w_matrix_reg_2__7__3_ ( .D(n2792), .CK(clk), .RN(rst_n), .Q(
        w_matrix[643]) );
  DFFRHQX1 w_matrix_reg_3__3__3_ ( .D(n2856), .CK(clk), .RN(rst_n), .Q(
        w_matrix[579]) );
  DFFRHQX1 w_matrix_reg_3__7__3_ ( .D(n2920), .CK(clk), .RN(rst_n), .Q(
        w_matrix[515]) );
  DFFRHQX1 w_matrix_reg_4__3__3_ ( .D(n2984), .CK(clk), .RN(rst_n), .Q(
        w_matrix[451]) );
  DFFRHQX1 w_matrix_reg_4__7__3_ ( .D(n3048), .CK(clk), .RN(rst_n), .Q(
        w_matrix[387]) );
  DFFRHQX1 w_matrix_reg_5__3__3_ ( .D(n3112), .CK(clk), .RN(rst_n), .Q(
        w_matrix[323]) );
  DFFRHQX1 w_matrix_reg_5__7__3_ ( .D(n3176), .CK(clk), .RN(rst_n), .Q(
        w_matrix[259]) );
  DFFRHQX1 w_matrix_reg_6__3__3_ ( .D(n3240), .CK(clk), .RN(rst_n), .Q(
        w_matrix[195]) );
  DFFRHQX1 w_matrix_reg_6__7__3_ ( .D(n3304), .CK(clk), .RN(rst_n), .Q(
        w_matrix[131]) );
  DFFRHQX1 w_matrix_reg_7__3__3_ ( .D(n3368), .CK(clk), .RN(rst_n), .Q(
        w_matrix[67]) );
  DFFRHQX1 w_matrix_reg_7__7__3_ ( .D(n3432), .CK(clk), .RN(rst_n), .Q(
        w_matrix[3]) );
  DFFRHQX1 w_matrix_reg_1__5__7_ ( .D(n2628), .CK(clk), .RN(rst_n), .Q(
        w_matrix[807]) );
  DFFRHQX1 w_matrix_reg_2__1__7_ ( .D(n2692), .CK(clk), .RN(rst_n), .Q(
        w_matrix[743]) );
  DFFRHQX1 w_matrix_reg_2__5__7_ ( .D(n2756), .CK(clk), .RN(rst_n), .Q(
        w_matrix[679]) );
  DFFRHQX1 w_matrix_reg_3__1__7_ ( .D(n2820), .CK(clk), .RN(rst_n), .Q(
        w_matrix[615]) );
  DFFRHQX1 w_matrix_reg_3__5__7_ ( .D(n2884), .CK(clk), .RN(rst_n), .Q(
        w_matrix[551]) );
  DFFRHQX1 w_matrix_reg_4__1__7_ ( .D(n2948), .CK(clk), .RN(rst_n), .Q(
        w_matrix[487]) );
  DFFRHQX1 w_matrix_reg_4__5__7_ ( .D(n3012), .CK(clk), .RN(rst_n), .Q(
        w_matrix[423]) );
  DFFRHQX1 w_matrix_reg_5__1__7_ ( .D(n3076), .CK(clk), .RN(rst_n), .Q(
        w_matrix[359]) );
  DFFRHQX1 w_matrix_reg_5__5__7_ ( .D(n3140), .CK(clk), .RN(rst_n), .Q(
        w_matrix[295]) );
  DFFRHQX1 w_matrix_reg_6__1__7_ ( .D(n3204), .CK(clk), .RN(rst_n), .Q(
        w_matrix[231]) );
  DFFRHQX1 w_matrix_reg_6__5__7_ ( .D(n3268), .CK(clk), .RN(rst_n), .Q(
        w_matrix[167]) );
  DFFRHQX1 w_matrix_reg_7__1__7_ ( .D(n3332), .CK(clk), .RN(rst_n), .Q(
        w_matrix[103]) );
  DFFRHQX1 w_matrix_reg_7__5__7_ ( .D(n3396), .CK(clk), .RN(rst_n), .Q(
        w_matrix[39]) );
  DFFRHQX1 w_matrix_reg_1__5__6_ ( .D(n2629), .CK(clk), .RN(rst_n), .Q(
        w_matrix[806]) );
  DFFRHQX1 w_matrix_reg_2__1__6_ ( .D(n2693), .CK(clk), .RN(rst_n), .Q(
        w_matrix[742]) );
  DFFRHQX1 w_matrix_reg_2__5__6_ ( .D(n2757), .CK(clk), .RN(rst_n), .Q(
        w_matrix[678]) );
  DFFRHQX1 w_matrix_reg_3__1__6_ ( .D(n2821), .CK(clk), .RN(rst_n), .Q(
        w_matrix[614]) );
  DFFRHQX1 w_matrix_reg_3__5__6_ ( .D(n2885), .CK(clk), .RN(rst_n), .Q(
        w_matrix[550]) );
  DFFRHQX1 w_matrix_reg_4__1__6_ ( .D(n2949), .CK(clk), .RN(rst_n), .Q(
        w_matrix[486]) );
  DFFRHQX1 w_matrix_reg_4__5__6_ ( .D(n3013), .CK(clk), .RN(rst_n), .Q(
        w_matrix[422]) );
  DFFRHQX1 w_matrix_reg_5__1__6_ ( .D(n3077), .CK(clk), .RN(rst_n), .Q(
        w_matrix[358]) );
  DFFRHQX1 w_matrix_reg_5__5__6_ ( .D(n3141), .CK(clk), .RN(rst_n), .Q(
        w_matrix[294]) );
  DFFRHQX1 w_matrix_reg_6__1__6_ ( .D(n3205), .CK(clk), .RN(rst_n), .Q(
        w_matrix[230]) );
  DFFRHQX1 w_matrix_reg_6__5__6_ ( .D(n3269), .CK(clk), .RN(rst_n), .Q(
        w_matrix[166]) );
  DFFRHQX1 w_matrix_reg_7__1__6_ ( .D(n3333), .CK(clk), .RN(rst_n), .Q(
        w_matrix[102]) );
  DFFRHQX1 w_matrix_reg_7__5__6_ ( .D(n3397), .CK(clk), .RN(rst_n), .Q(
        w_matrix[38]) );
  DFFRHQX1 w_matrix_reg_1__5__5_ ( .D(n2630), .CK(clk), .RN(rst_n), .Q(
        w_matrix[805]) );
  DFFRHQX1 w_matrix_reg_2__1__5_ ( .D(n2694), .CK(clk), .RN(rst_n), .Q(
        w_matrix[741]) );
  DFFRHQX1 w_matrix_reg_2__5__5_ ( .D(n2758), .CK(clk), .RN(rst_n), .Q(
        w_matrix[677]) );
  DFFRHQX1 w_matrix_reg_3__1__5_ ( .D(n2822), .CK(clk), .RN(rst_n), .Q(
        w_matrix[613]) );
  DFFRHQX1 w_matrix_reg_3__5__5_ ( .D(n2886), .CK(clk), .RN(rst_n), .Q(
        w_matrix[549]) );
  DFFRHQX1 w_matrix_reg_4__1__5_ ( .D(n2950), .CK(clk), .RN(rst_n), .Q(
        w_matrix[485]) );
  DFFRHQX1 w_matrix_reg_4__5__5_ ( .D(n3014), .CK(clk), .RN(rst_n), .Q(
        w_matrix[421]) );
  DFFRHQX1 w_matrix_reg_5__1__5_ ( .D(n3078), .CK(clk), .RN(rst_n), .Q(
        w_matrix[357]) );
  DFFRHQX1 w_matrix_reg_5__5__5_ ( .D(n3142), .CK(clk), .RN(rst_n), .Q(
        w_matrix[293]) );
  DFFRHQX1 w_matrix_reg_6__1__5_ ( .D(n3206), .CK(clk), .RN(rst_n), .Q(
        w_matrix[229]) );
  DFFRHQX1 w_matrix_reg_6__5__5_ ( .D(n3270), .CK(clk), .RN(rst_n), .Q(
        w_matrix[165]) );
  DFFRHQX1 w_matrix_reg_7__1__5_ ( .D(n3334), .CK(clk), .RN(rst_n), .Q(
        w_matrix[101]) );
  DFFRHQX1 w_matrix_reg_7__5__5_ ( .D(n3398), .CK(clk), .RN(rst_n), .Q(
        w_matrix[37]) );
  DFFRHQX1 w_matrix_reg_1__5__4_ ( .D(n2631), .CK(clk), .RN(rst_n), .Q(
        w_matrix[804]) );
  DFFRHQX1 w_matrix_reg_2__1__4_ ( .D(n2695), .CK(clk), .RN(rst_n), .Q(
        w_matrix[740]) );
  DFFRHQX1 w_matrix_reg_2__5__4_ ( .D(n2759), .CK(clk), .RN(rst_n), .Q(
        w_matrix[676]) );
  DFFRHQX1 w_matrix_reg_3__1__4_ ( .D(n2823), .CK(clk), .RN(rst_n), .Q(
        w_matrix[612]) );
  DFFRHQX1 w_matrix_reg_3__5__4_ ( .D(n2887), .CK(clk), .RN(rst_n), .Q(
        w_matrix[548]) );
  DFFRHQX1 w_matrix_reg_4__1__4_ ( .D(n2951), .CK(clk), .RN(rst_n), .Q(
        w_matrix[484]) );
  DFFRHQX1 w_matrix_reg_4__5__4_ ( .D(n3015), .CK(clk), .RN(rst_n), .Q(
        w_matrix[420]) );
  DFFRHQX1 w_matrix_reg_5__1__4_ ( .D(n3079), .CK(clk), .RN(rst_n), .Q(
        w_matrix[356]) );
  DFFRHQX1 w_matrix_reg_5__5__4_ ( .D(n3143), .CK(clk), .RN(rst_n), .Q(
        w_matrix[292]) );
  DFFRHQX1 w_matrix_reg_6__1__4_ ( .D(n3207), .CK(clk), .RN(rst_n), .Q(
        w_matrix[228]) );
  DFFRHQX1 w_matrix_reg_6__5__4_ ( .D(n3271), .CK(clk), .RN(rst_n), .Q(
        w_matrix[164]) );
  DFFRHQX1 w_matrix_reg_7__1__4_ ( .D(n3335), .CK(clk), .RN(rst_n), .Q(
        w_matrix[100]) );
  DFFRHQX1 w_matrix_reg_7__5__4_ ( .D(n3399), .CK(clk), .RN(rst_n), .Q(
        w_matrix[36]) );
  DFFRHQX1 w_matrix_reg_1__5__3_ ( .D(n2632), .CK(clk), .RN(rst_n), .Q(
        w_matrix[803]) );
  DFFRHQX1 w_matrix_reg_2__1__3_ ( .D(n2696), .CK(clk), .RN(rst_n), .Q(
        w_matrix[739]) );
  DFFRHQX1 w_matrix_reg_2__5__3_ ( .D(n2760), .CK(clk), .RN(rst_n), .Q(
        w_matrix[675]) );
  DFFRHQX1 w_matrix_reg_3__1__3_ ( .D(n2824), .CK(clk), .RN(rst_n), .Q(
        w_matrix[611]) );
  DFFRHQX1 w_matrix_reg_3__5__3_ ( .D(n2888), .CK(clk), .RN(rst_n), .Q(
        w_matrix[547]) );
  DFFRHQX1 w_matrix_reg_4__1__3_ ( .D(n2952), .CK(clk), .RN(rst_n), .Q(
        w_matrix[483]) );
  DFFRHQX1 w_matrix_reg_4__5__3_ ( .D(n3016), .CK(clk), .RN(rst_n), .Q(
        w_matrix[419]) );
  DFFRHQX1 w_matrix_reg_5__1__3_ ( .D(n3080), .CK(clk), .RN(rst_n), .Q(
        w_matrix[355]) );
  DFFRHQX1 w_matrix_reg_5__5__3_ ( .D(n3144), .CK(clk), .RN(rst_n), .Q(
        w_matrix[291]) );
  DFFRHQX1 w_matrix_reg_6__1__3_ ( .D(n3208), .CK(clk), .RN(rst_n), .Q(
        w_matrix[227]) );
  DFFRHQX1 w_matrix_reg_6__5__3_ ( .D(n3272), .CK(clk), .RN(rst_n), .Q(
        w_matrix[163]) );
  DFFRHQX1 w_matrix_reg_7__1__3_ ( .D(n3336), .CK(clk), .RN(rst_n), .Q(
        w_matrix[99]) );
  DFFRHQX1 w_matrix_reg_7__5__3_ ( .D(n3400), .CK(clk), .RN(rst_n), .Q(
        w_matrix[35]) );
  DFFRHQX1 w_matrix_reg_1__5__2_ ( .D(n2633), .CK(clk), .RN(rst_n), .Q(
        w_matrix[802]) );
  DFFRHQX1 w_matrix_reg_2__1__2_ ( .D(n2697), .CK(clk), .RN(rst_n), .Q(
        w_matrix[738]) );
  DFFRHQX1 w_matrix_reg_2__5__2_ ( .D(n2761), .CK(clk), .RN(rst_n), .Q(
        w_matrix[674]) );
  DFFRHQX1 w_matrix_reg_3__1__2_ ( .D(n2825), .CK(clk), .RN(rst_n), .Q(
        w_matrix[610]) );
  DFFRHQX1 w_matrix_reg_3__5__2_ ( .D(n2889), .CK(clk), .RN(rst_n), .Q(
        w_matrix[546]) );
  DFFRHQX1 w_matrix_reg_4__1__2_ ( .D(n2953), .CK(clk), .RN(rst_n), .Q(
        w_matrix[482]) );
  DFFRHQX1 w_matrix_reg_4__5__2_ ( .D(n3017), .CK(clk), .RN(rst_n), .Q(
        w_matrix[418]) );
  DFFRHQX1 w_matrix_reg_5__1__2_ ( .D(n3081), .CK(clk), .RN(rst_n), .Q(
        w_matrix[354]) );
  DFFRHQX1 w_matrix_reg_5__5__2_ ( .D(n3145), .CK(clk), .RN(rst_n), .Q(
        w_matrix[290]) );
  DFFRHQX1 w_matrix_reg_6__1__2_ ( .D(n3209), .CK(clk), .RN(rst_n), .Q(
        w_matrix[226]) );
  DFFRHQX1 w_matrix_reg_6__5__2_ ( .D(n3273), .CK(clk), .RN(rst_n), .Q(
        w_matrix[162]) );
  DFFRHQX1 w_matrix_reg_7__1__2_ ( .D(n3337), .CK(clk), .RN(rst_n), .Q(
        w_matrix[98]) );
  DFFRHQX1 w_matrix_reg_7__5__2_ ( .D(n3401), .CK(clk), .RN(rst_n), .Q(
        w_matrix[34]) );
  DFFRHQX1 w_matrix_reg_1__5__1_ ( .D(n2634), .CK(clk), .RN(rst_n), .Q(
        w_matrix[801]) );
  DFFRHQX1 w_matrix_reg_2__1__1_ ( .D(n2698), .CK(clk), .RN(rst_n), .Q(
        w_matrix[737]) );
  DFFRHQX1 w_matrix_reg_2__5__1_ ( .D(n2762), .CK(clk), .RN(rst_n), .Q(
        w_matrix[673]) );
  DFFRHQX1 w_matrix_reg_3__1__1_ ( .D(n2826), .CK(clk), .RN(rst_n), .Q(
        w_matrix[609]) );
  DFFRHQX1 w_matrix_reg_3__5__1_ ( .D(n2890), .CK(clk), .RN(rst_n), .Q(
        w_matrix[545]) );
  DFFRHQX1 w_matrix_reg_4__1__1_ ( .D(n2954), .CK(clk), .RN(rst_n), .Q(
        w_matrix[481]) );
  DFFRHQX1 w_matrix_reg_4__5__1_ ( .D(n3018), .CK(clk), .RN(rst_n), .Q(
        w_matrix[417]) );
  DFFRHQX1 w_matrix_reg_5__1__1_ ( .D(n3082), .CK(clk), .RN(rst_n), .Q(
        w_matrix[353]) );
  DFFRHQX1 w_matrix_reg_5__5__1_ ( .D(n3146), .CK(clk), .RN(rst_n), .Q(
        w_matrix[289]) );
  DFFRHQX1 w_matrix_reg_6__1__1_ ( .D(n3210), .CK(clk), .RN(rst_n), .Q(
        w_matrix[225]) );
  DFFRHQX1 w_matrix_reg_6__5__1_ ( .D(n3274), .CK(clk), .RN(rst_n), .Q(
        w_matrix[161]) );
  DFFRHQX1 w_matrix_reg_7__1__1_ ( .D(n3338), .CK(clk), .RN(rst_n), .Q(
        w_matrix[97]) );
  DFFRHQX1 w_matrix_reg_7__5__1_ ( .D(n3402), .CK(clk), .RN(rst_n), .Q(
        w_matrix[33]) );
  DFFRHQX1 w_matrix_reg_1__3__2_ ( .D(n2601), .CK(clk), .RN(rst_n), .Q(
        w_matrix[834]) );
  DFFRHQX1 w_matrix_reg_1__7__2_ ( .D(n2665), .CK(clk), .RN(rst_n), .Q(
        w_matrix[770]) );
  DFFRHQX1 w_matrix_reg_2__3__2_ ( .D(n2729), .CK(clk), .RN(rst_n), .Q(
        w_matrix[706]) );
  DFFRHQX1 w_matrix_reg_2__7__2_ ( .D(n2793), .CK(clk), .RN(rst_n), .Q(
        w_matrix[642]) );
  DFFRHQX1 w_matrix_reg_3__3__2_ ( .D(n2857), .CK(clk), .RN(rst_n), .Q(
        w_matrix[578]) );
  DFFRHQX1 w_matrix_reg_3__7__2_ ( .D(n2921), .CK(clk), .RN(rst_n), .Q(
        w_matrix[514]) );
  DFFRHQX1 w_matrix_reg_4__3__2_ ( .D(n2985), .CK(clk), .RN(rst_n), .Q(
        w_matrix[450]) );
  DFFRHQX1 w_matrix_reg_4__7__2_ ( .D(n3049), .CK(clk), .RN(rst_n), .Q(
        w_matrix[386]) );
  DFFRHQX1 w_matrix_reg_5__3__2_ ( .D(n3113), .CK(clk), .RN(rst_n), .Q(
        w_matrix[322]) );
  DFFRHQX1 w_matrix_reg_5__7__2_ ( .D(n3177), .CK(clk), .RN(rst_n), .Q(
        w_matrix[258]) );
  DFFRHQX1 w_matrix_reg_6__3__2_ ( .D(n3241), .CK(clk), .RN(rst_n), .Q(
        w_matrix[194]) );
  DFFRHQX1 w_matrix_reg_6__7__2_ ( .D(n3305), .CK(clk), .RN(rst_n), .Q(
        w_matrix[130]) );
  DFFRHQX1 w_matrix_reg_7__3__2_ ( .D(n3369), .CK(clk), .RN(rst_n), .Q(
        w_matrix[66]) );
  DFFRHQX1 w_matrix_reg_7__7__2_ ( .D(n3433), .CK(clk), .RN(rst_n), .Q(
        w_matrix[2]) );
  DFFRHQX1 w_matrix_reg_1__2__7_ ( .D(n2580), .CK(clk), .RN(rst_n), .Q(
        w_matrix[855]) );
  DFFRHQX1 w_matrix_reg_1__6__7_ ( .D(n2644), .CK(clk), .RN(rst_n), .Q(
        w_matrix[791]) );
  DFFRHQX1 w_matrix_reg_2__2__7_ ( .D(n2708), .CK(clk), .RN(rst_n), .Q(
        w_matrix[727]) );
  DFFRHQX1 w_matrix_reg_2__6__7_ ( .D(n2772), .CK(clk), .RN(rst_n), .Q(
        w_matrix[663]) );
  DFFRHQX1 w_matrix_reg_3__2__7_ ( .D(n2836), .CK(clk), .RN(rst_n), .Q(
        w_matrix[599]) );
  DFFRHQX1 w_matrix_reg_3__6__7_ ( .D(n2900), .CK(clk), .RN(rst_n), .Q(
        w_matrix[535]) );
  DFFRHQX1 w_matrix_reg_4__2__7_ ( .D(n2964), .CK(clk), .RN(rst_n), .Q(
        w_matrix[471]) );
  DFFRHQX1 w_matrix_reg_4__6__7_ ( .D(n3028), .CK(clk), .RN(rst_n), .Q(
        w_matrix[407]) );
  DFFRHQX1 w_matrix_reg_5__2__7_ ( .D(n3092), .CK(clk), .RN(rst_n), .Q(
        w_matrix[343]) );
  DFFRHQX1 w_matrix_reg_5__6__7_ ( .D(n3156), .CK(clk), .RN(rst_n), .Q(
        w_matrix[279]) );
  DFFRHQX1 w_matrix_reg_6__2__7_ ( .D(n3220), .CK(clk), .RN(rst_n), .Q(
        w_matrix[215]) );
  DFFRHQX1 w_matrix_reg_6__6__7_ ( .D(n3284), .CK(clk), .RN(rst_n), .Q(
        w_matrix[151]) );
  DFFRHQX1 w_matrix_reg_7__2__7_ ( .D(n3348), .CK(clk), .RN(rst_n), .Q(
        w_matrix[87]) );
  DFFRHQX1 w_matrix_reg_7__6__7_ ( .D(n3412), .CK(clk), .RN(rst_n), .Q(
        w_matrix[23]) );
  DFFRHQX1 w_matrix_reg_1__2__6_ ( .D(n2581), .CK(clk), .RN(rst_n), .Q(
        w_matrix[854]) );
  DFFRHQX1 w_matrix_reg_1__6__6_ ( .D(n2645), .CK(clk), .RN(rst_n), .Q(
        w_matrix[790]) );
  DFFRHQX1 w_matrix_reg_2__2__6_ ( .D(n2709), .CK(clk), .RN(rst_n), .Q(
        w_matrix[726]) );
  DFFRHQX1 w_matrix_reg_2__6__6_ ( .D(n2773), .CK(clk), .RN(rst_n), .Q(
        w_matrix[662]) );
  DFFRHQX1 w_matrix_reg_3__2__6_ ( .D(n2837), .CK(clk), .RN(rst_n), .Q(
        w_matrix[598]) );
  DFFRHQX1 w_matrix_reg_3__6__6_ ( .D(n2901), .CK(clk), .RN(rst_n), .Q(
        w_matrix[534]) );
  DFFRHQX1 w_matrix_reg_4__2__6_ ( .D(n2965), .CK(clk), .RN(rst_n), .Q(
        w_matrix[470]) );
  DFFRHQX1 w_matrix_reg_4__6__6_ ( .D(n3029), .CK(clk), .RN(rst_n), .Q(
        w_matrix[406]) );
  DFFRHQX1 w_matrix_reg_5__2__6_ ( .D(n3093), .CK(clk), .RN(rst_n), .Q(
        w_matrix[342]) );
  DFFRHQX1 w_matrix_reg_5__6__6_ ( .D(n3157), .CK(clk), .RN(rst_n), .Q(
        w_matrix[278]) );
  DFFRHQX1 w_matrix_reg_6__2__6_ ( .D(n3221), .CK(clk), .RN(rst_n), .Q(
        w_matrix[214]) );
  DFFRHQX1 w_matrix_reg_6__6__6_ ( .D(n3285), .CK(clk), .RN(rst_n), .Q(
        w_matrix[150]) );
  DFFRHQX1 w_matrix_reg_7__2__6_ ( .D(n3349), .CK(clk), .RN(rst_n), .Q(
        w_matrix[86]) );
  DFFRHQX1 w_matrix_reg_7__6__6_ ( .D(n3413), .CK(clk), .RN(rst_n), .Q(
        w_matrix[22]) );
  DFFRHQX1 w_matrix_reg_1__2__5_ ( .D(n2582), .CK(clk), .RN(rst_n), .Q(
        w_matrix[853]) );
  DFFRHQX1 w_matrix_reg_1__6__5_ ( .D(n2646), .CK(clk), .RN(rst_n), .Q(
        w_matrix[789]) );
  DFFRHQX1 w_matrix_reg_2__2__5_ ( .D(n2710), .CK(clk), .RN(rst_n), .Q(
        w_matrix[725]) );
  DFFRHQX1 w_matrix_reg_2__6__5_ ( .D(n2774), .CK(clk), .RN(rst_n), .Q(
        w_matrix[661]) );
  DFFRHQX1 w_matrix_reg_3__2__5_ ( .D(n2838), .CK(clk), .RN(rst_n), .Q(
        w_matrix[597]) );
  DFFRHQX1 w_matrix_reg_3__6__5_ ( .D(n2902), .CK(clk), .RN(rst_n), .Q(
        w_matrix[533]) );
  DFFRHQX1 w_matrix_reg_4__2__5_ ( .D(n2966), .CK(clk), .RN(rst_n), .Q(
        w_matrix[469]) );
  DFFRHQX1 w_matrix_reg_4__6__5_ ( .D(n3030), .CK(clk), .RN(rst_n), .Q(
        w_matrix[405]) );
  DFFRHQX1 w_matrix_reg_5__2__5_ ( .D(n3094), .CK(clk), .RN(rst_n), .Q(
        w_matrix[341]) );
  DFFRHQX1 w_matrix_reg_5__6__5_ ( .D(n3158), .CK(clk), .RN(rst_n), .Q(
        w_matrix[277]) );
  DFFRHQX1 w_matrix_reg_6__2__5_ ( .D(n3222), .CK(clk), .RN(rst_n), .Q(
        w_matrix[213]) );
  DFFRHQX1 w_matrix_reg_6__6__5_ ( .D(n3286), .CK(clk), .RN(rst_n), .Q(
        w_matrix[149]) );
  DFFRHQX1 w_matrix_reg_7__2__5_ ( .D(n3350), .CK(clk), .RN(rst_n), .Q(
        w_matrix[85]) );
  DFFRHQX1 w_matrix_reg_7__6__5_ ( .D(n3414), .CK(clk), .RN(rst_n), .Q(
        w_matrix[21]) );
  DFFRHQX1 w_matrix_reg_1__2__4_ ( .D(n2583), .CK(clk), .RN(rst_n), .Q(
        w_matrix[852]) );
  DFFRHQX1 w_matrix_reg_1__6__4_ ( .D(n2647), .CK(clk), .RN(rst_n), .Q(
        w_matrix[788]) );
  DFFRHQX1 w_matrix_reg_2__2__4_ ( .D(n2711), .CK(clk), .RN(rst_n), .Q(
        w_matrix[724]) );
  DFFRHQX1 w_matrix_reg_2__6__4_ ( .D(n2775), .CK(clk), .RN(rst_n), .Q(
        w_matrix[660]) );
  DFFRHQX1 w_matrix_reg_3__2__4_ ( .D(n2839), .CK(clk), .RN(rst_n), .Q(
        w_matrix[596]) );
  DFFRHQX1 w_matrix_reg_3__6__4_ ( .D(n2903), .CK(clk), .RN(rst_n), .Q(
        w_matrix[532]) );
  DFFRHQX1 w_matrix_reg_4__2__4_ ( .D(n2967), .CK(clk), .RN(rst_n), .Q(
        w_matrix[468]) );
  DFFRHQX1 w_matrix_reg_4__6__4_ ( .D(n3031), .CK(clk), .RN(rst_n), .Q(
        w_matrix[404]) );
  DFFRHQX1 w_matrix_reg_5__2__4_ ( .D(n3095), .CK(clk), .RN(rst_n), .Q(
        w_matrix[340]) );
  DFFRHQX1 w_matrix_reg_5__6__4_ ( .D(n3159), .CK(clk), .RN(rst_n), .Q(
        w_matrix[276]) );
  DFFRHQX1 w_matrix_reg_6__2__4_ ( .D(n3223), .CK(clk), .RN(rst_n), .Q(
        w_matrix[212]) );
  DFFRHQX1 w_matrix_reg_6__6__4_ ( .D(n3287), .CK(clk), .RN(rst_n), .Q(
        w_matrix[148]) );
  DFFRHQX1 w_matrix_reg_7__2__4_ ( .D(n3351), .CK(clk), .RN(rst_n), .Q(
        w_matrix[84]) );
  DFFRHQX1 w_matrix_reg_7__6__4_ ( .D(n3415), .CK(clk), .RN(rst_n), .Q(
        w_matrix[20]) );
  DFFRHQX1 w_matrix_reg_1__3__1_ ( .D(n2602), .CK(clk), .RN(rst_n), .Q(
        w_matrix[833]) );
  DFFRHQX1 w_matrix_reg_1__7__1_ ( .D(n2666), .CK(clk), .RN(rst_n), .Q(
        w_matrix[769]) );
  DFFRHQX1 w_matrix_reg_2__3__1_ ( .D(n2730), .CK(clk), .RN(rst_n), .Q(
        w_matrix[705]) );
  DFFRHQX1 w_matrix_reg_2__7__1_ ( .D(n2794), .CK(clk), .RN(rst_n), .Q(
        w_matrix[641]) );
  DFFRHQX1 w_matrix_reg_3__3__1_ ( .D(n2858), .CK(clk), .RN(rst_n), .Q(
        w_matrix[577]) );
  DFFRHQX1 w_matrix_reg_3__7__1_ ( .D(n2922), .CK(clk), .RN(rst_n), .Q(
        w_matrix[513]) );
  DFFRHQX1 w_matrix_reg_4__3__1_ ( .D(n2986), .CK(clk), .RN(rst_n), .Q(
        w_matrix[449]) );
  DFFRHQX1 w_matrix_reg_4__7__1_ ( .D(n3050), .CK(clk), .RN(rst_n), .Q(
        w_matrix[385]) );
  DFFRHQX1 w_matrix_reg_5__3__1_ ( .D(n3114), .CK(clk), .RN(rst_n), .Q(
        w_matrix[321]) );
  DFFRHQX1 w_matrix_reg_5__7__1_ ( .D(n3178), .CK(clk), .RN(rst_n), .Q(
        w_matrix[257]) );
  DFFRHQX1 w_matrix_reg_6__3__1_ ( .D(n3242), .CK(clk), .RN(rst_n), .Q(
        w_matrix[193]) );
  DFFRHQX1 w_matrix_reg_6__7__1_ ( .D(n3306), .CK(clk), .RN(rst_n), .Q(
        w_matrix[129]) );
  DFFRHQX1 w_matrix_reg_7__3__1_ ( .D(n3370), .CK(clk), .RN(rst_n), .Q(
        w_matrix[65]) );
  DFFRHQX1 w_matrix_reg_7__7__1_ ( .D(n3434), .CK(clk), .RN(rst_n), .Q(
        w_matrix[1]) );
  DFFRHQX1 w_matrix_reg_1__2__3_ ( .D(n2584), .CK(clk), .RN(rst_n), .Q(
        w_matrix[851]) );
  DFFRHQX1 w_matrix_reg_1__6__3_ ( .D(n2648), .CK(clk), .RN(rst_n), .Q(
        w_matrix[787]) );
  DFFRHQX1 w_matrix_reg_2__2__3_ ( .D(n2712), .CK(clk), .RN(rst_n), .Q(
        w_matrix[723]) );
  DFFRHQX1 w_matrix_reg_2__6__3_ ( .D(n2776), .CK(clk), .RN(rst_n), .Q(
        w_matrix[659]) );
  DFFRHQX1 w_matrix_reg_3__2__3_ ( .D(n2840), .CK(clk), .RN(rst_n), .Q(
        w_matrix[595]) );
  DFFRHQX1 w_matrix_reg_3__6__3_ ( .D(n2904), .CK(clk), .RN(rst_n), .Q(
        w_matrix[531]) );
  DFFRHQX1 w_matrix_reg_4__2__3_ ( .D(n2968), .CK(clk), .RN(rst_n), .Q(
        w_matrix[467]) );
  DFFRHQX1 w_matrix_reg_4__6__3_ ( .D(n3032), .CK(clk), .RN(rst_n), .Q(
        w_matrix[403]) );
  DFFRHQX1 w_matrix_reg_5__2__3_ ( .D(n3096), .CK(clk), .RN(rst_n), .Q(
        w_matrix[339]) );
  DFFRHQX1 w_matrix_reg_5__6__3_ ( .D(n3160), .CK(clk), .RN(rst_n), .Q(
        w_matrix[275]) );
  DFFRHQX1 w_matrix_reg_6__2__3_ ( .D(n3224), .CK(clk), .RN(rst_n), .Q(
        w_matrix[211]) );
  DFFRHQX1 w_matrix_reg_6__6__3_ ( .D(n3288), .CK(clk), .RN(rst_n), .Q(
        w_matrix[147]) );
  DFFRHQX1 w_matrix_reg_7__2__3_ ( .D(n3352), .CK(clk), .RN(rst_n), .Q(
        w_matrix[83]) );
  DFFRHQX1 w_matrix_reg_7__6__3_ ( .D(n3416), .CK(clk), .RN(rst_n), .Q(
        w_matrix[19]) );
  DFFRHQX1 w_matrix_reg_1__2__2_ ( .D(n2585), .CK(clk), .RN(rst_n), .Q(
        w_matrix[850]) );
  DFFRHQX1 w_matrix_reg_1__6__2_ ( .D(n2649), .CK(clk), .RN(rst_n), .Q(
        w_matrix[786]) );
  DFFRHQX1 w_matrix_reg_2__2__2_ ( .D(n2713), .CK(clk), .RN(rst_n), .Q(
        w_matrix[722]) );
  DFFRHQX1 w_matrix_reg_2__6__2_ ( .D(n2777), .CK(clk), .RN(rst_n), .Q(
        w_matrix[658]) );
  DFFRHQX1 w_matrix_reg_3__2__2_ ( .D(n2841), .CK(clk), .RN(rst_n), .Q(
        w_matrix[594]) );
  DFFRHQX1 w_matrix_reg_3__6__2_ ( .D(n2905), .CK(clk), .RN(rst_n), .Q(
        w_matrix[530]) );
  DFFRHQX1 w_matrix_reg_4__2__2_ ( .D(n2969), .CK(clk), .RN(rst_n), .Q(
        w_matrix[466]) );
  DFFRHQX1 w_matrix_reg_4__6__2_ ( .D(n3033), .CK(clk), .RN(rst_n), .Q(
        w_matrix[402]) );
  DFFRHQX1 w_matrix_reg_5__2__2_ ( .D(n3097), .CK(clk), .RN(rst_n), .Q(
        w_matrix[338]) );
  DFFRHQX1 w_matrix_reg_5__6__2_ ( .D(n3161), .CK(clk), .RN(rst_n), .Q(
        w_matrix[274]) );
  DFFRHQX1 w_matrix_reg_6__2__2_ ( .D(n3225), .CK(clk), .RN(rst_n), .Q(
        w_matrix[210]) );
  DFFRHQX1 w_matrix_reg_6__6__2_ ( .D(n3289), .CK(clk), .RN(rst_n), .Q(
        w_matrix[146]) );
  DFFRHQX1 w_matrix_reg_7__2__2_ ( .D(n3353), .CK(clk), .RN(rst_n), .Q(
        w_matrix[82]) );
  DFFRHQX1 w_matrix_reg_7__6__2_ ( .D(n3417), .CK(clk), .RN(rst_n), .Q(
        w_matrix[18]) );
  DFFRHQX1 w_matrix_reg_1__2__1_ ( .D(n2586), .CK(clk), .RN(rst_n), .Q(
        w_matrix[849]) );
  DFFRHQX1 w_matrix_reg_1__6__1_ ( .D(n2650), .CK(clk), .RN(rst_n), .Q(
        w_matrix[785]) );
  DFFRHQX1 w_matrix_reg_2__2__1_ ( .D(n2714), .CK(clk), .RN(rst_n), .Q(
        w_matrix[721]) );
  DFFRHQX1 w_matrix_reg_2__6__1_ ( .D(n2778), .CK(clk), .RN(rst_n), .Q(
        w_matrix[657]) );
  DFFRHQX1 w_matrix_reg_3__2__1_ ( .D(n2842), .CK(clk), .RN(rst_n), .Q(
        w_matrix[593]) );
  DFFRHQX1 w_matrix_reg_3__6__1_ ( .D(n2906), .CK(clk), .RN(rst_n), .Q(
        w_matrix[529]) );
  DFFRHQX1 w_matrix_reg_4__2__1_ ( .D(n2970), .CK(clk), .RN(rst_n), .Q(
        w_matrix[465]) );
  DFFRHQX1 w_matrix_reg_4__6__1_ ( .D(n3034), .CK(clk), .RN(rst_n), .Q(
        w_matrix[401]) );
  DFFRHQX1 w_matrix_reg_5__2__1_ ( .D(n3098), .CK(clk), .RN(rst_n), .Q(
        w_matrix[337]) );
  DFFRHQX1 w_matrix_reg_5__6__1_ ( .D(n3162), .CK(clk), .RN(rst_n), .Q(
        w_matrix[273]) );
  DFFRHQX1 w_matrix_reg_6__2__1_ ( .D(n3226), .CK(clk), .RN(rst_n), .Q(
        w_matrix[209]) );
  DFFRHQX1 w_matrix_reg_6__6__1_ ( .D(n3290), .CK(clk), .RN(rst_n), .Q(
        w_matrix[145]) );
  DFFRHQX1 w_matrix_reg_7__2__1_ ( .D(n3354), .CK(clk), .RN(rst_n), .Q(
        w_matrix[81]) );
  DFFRHQX1 w_matrix_reg_7__6__1_ ( .D(n3418), .CK(clk), .RN(rst_n), .Q(
        w_matrix[17]) );
  DFFRHQX1 inA51_reg_0_ ( .D(N11773), .CK(clk), .RN(rst_n), .Q(inA51[0]) );
  DFFRHQX1 inA61_reg_0_ ( .D(N11870), .CK(clk), .RN(rst_n), .Q(inA61[0]) );
  DFFRHQX1 inA31_reg_0_ ( .D(N11584), .CK(clk), .RN(rst_n), .Q(inA31[0]) );
  DFFRHQX1 inA71_reg_0_ ( .D(N11964), .CK(clk), .RN(rst_n), .Q(inA71[0]) );
  DFFRHQX1 inA21_reg_0_ ( .D(N11490), .CK(clk), .RN(rst_n), .Q(inA21[0]) );
  DFFRHQX1 inA41_reg_0_ ( .D(N11681), .CK(clk), .RN(rst_n), .Q(inA41[0]) );
  DFFRHQX1 inA81_reg_0_ ( .D(N12060), .CK(clk), .RN(rst_n), .Q(inA81[0]) );
  DFFRHQX1 w_matrix_reg_1__0__0_ ( .D(n2555), .CK(clk), .RN(rst_n), .Q(
        w_matrix[880]) );
  DFFRX2 w_matrix_reg_1__1__0_ ( .D(n2571), .CK(clk), .RN(rst_n), .Q(
        w_matrix[864]), .QN(n673) );
  DFFRHQX1 inA51_reg_1_ ( .D(N11774), .CK(clk), .RN(rst_n), .Q(inA51[1]) );
  DFFRHQX1 inA61_reg_1_ ( .D(N11871), .CK(clk), .RN(rst_n), .Q(inA61[1]) );
  DFFRHQX1 inA21_reg_1_ ( .D(N11491), .CK(clk), .RN(rst_n), .Q(inA21[1]) );
  DFFRHQX1 inA41_reg_1_ ( .D(N11682), .CK(clk), .RN(rst_n), .Q(inA41[1]) );
  DFFRHQX1 inA81_reg_1_ ( .D(N12061), .CK(clk), .RN(rst_n), .Q(inA81[1]) );
  DFFRHQX1 inA31_reg_1_ ( .D(N11585), .CK(clk), .RN(rst_n), .Q(inA31[1]) );
  DFFRHQX1 inA71_reg_1_ ( .D(N11965), .CK(clk), .RN(rst_n), .Q(inA71[1]) );
  DFFRHQX1 in_64_reg_63_ ( .D(N1225), .CK(clk), .RN(rst_n), .Q(in_64[63]) );
  DFFRHQX1 in_matrix_cnt_reg_0_ ( .D(n5792), .CK(clk), .RN(rst_n), .Q(
        in_matrix_cnt[0]) );
  DFFRHQX1 in_matrix_cnt_reg_1_ ( .D(n5793), .CK(clk), .RN(rst_n), .Q(
        in_matrix_cnt[1]) );
  DFFRHQX1 in_matrix_cnt_reg_2_ ( .D(n5794), .CK(clk), .RN(rst_n), .Q(
        in_matrix_cnt[2]) );
  DFFRHQX1 in_matrix_cnt_reg_3_ ( .D(n5795), .CK(clk), .RN(rst_n), .Q(
        in_matrix_cnt[3]) );
  DFFRHQX1 calweight_addr_reg_0_ ( .D(n5812), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[0]) );
  DFFRHQX1 calin_addr_reg_0_ ( .D(n5803), .CK(clk), .RN(rst_n), .Q(
        calin_addr[0]) );
  DFFSX1 in_addr_cnt_reg_4_ ( .D(n4465), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[4]) );
  DFFSX1 in_addr_cnt_reg_5_ ( .D(n4464), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[5]) );
  DFFSX1 in_addr_cnt_reg_7_ ( .D(n4462), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[7]) );
  DFFSX1 in_addr_cnt_reg_6_ ( .D(n4463), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[6]) );
  DFFSX1 in_addr_cnt_reg_3_ ( .D(n4466), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[3]) );
  DFFSX1 in_addr_cnt_reg_2_ ( .D(n4467), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[2]) );
  DFFRHQX1 in_cnt_reg_0_ ( .D(n5831), .CK(clk), .RN(rst_n), .Q(in_cnt[0]) );
  DFFRHQX1 in_cnt_reg_1_ ( .D(n5830), .CK(clk), .RN(rst_n), .Q(in_cnt[1]) );
  DFFRHQX1 in_cnt_reg_2_ ( .D(n5829), .CK(clk), .RN(rst_n), .Q(in_cnt[2]) );
  DFFRHQX1 in_cnt_reg_3_ ( .D(n5828), .CK(clk), .RN(rst_n), .Q(in_cnt[3]) );
  DFFRHQX1 in_cnt_64_reg_0_ ( .D(N1040), .CK(clk), .RN(rst_n), .Q(in_cnt_64[0]) );
  DFFRHQX1 in_cnt_64_reg_4_ ( .D(N1044), .CK(clk), .RN(rst_n), .Q(in_cnt_64[4]) );
  DFFRHQX1 in_cnt_reg_5_ ( .D(n5826), .CK(clk), .RN(rst_n), .Q(in_cnt[5]) );
  DFFRHQX1 in_cnt_reg_6_ ( .D(n5825), .CK(clk), .RN(rst_n), .Q(in_cnt[6]) );
  DFFRHQX1 in_cnt_reg_4_ ( .D(n5827), .CK(clk), .RN(rst_n), .Q(in_cnt[4]) );
  DFFRHQX1 in_cnt_64_reg_3_ ( .D(N1043), .CK(clk), .RN(rst_n), .Q(in_cnt_64[3]) );
  DFFRHQX1 in_cnt_64_reg_1_ ( .D(N1041), .CK(clk), .RN(rst_n), .Q(in_cnt_64[1]) );
  DFFRHQX1 in_cnt_64_reg_2_ ( .D(N1042), .CK(clk), .RN(rst_n), .Q(in_cnt_64[2]) );
  DFFSX1 in_addr_cnt_reg_0_ ( .D(n4469), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[0]) );
  DFFSX1 in_addr_cnt_reg_1_ ( .D(n4468), .CK(clk), .SN(rst_n), .Q(
        in_addr_cnt[1]) );
  DFFRHQX1 store_cnt_reg_3_ ( .D(N14273), .CK(clk), .RN(rst_n), .Q(
        store_cnt[3]) );
  DFFRHQX1 outset_cnt_reg_0_ ( .D(n4472), .CK(clk), .RN(rst_n), .Q(N942) );
  DFFRHQX1 m_size_reg_0_ ( .D(n4470), .CK(clk), .RN(rst_n), .Q(m_size[0]) );
  DFFRHQX1 out_cnt_reg_0_ ( .D(n5839), .CK(clk), .RN(rst_n), .Q(out_cnt[0]) );
  DFFRHQX1 cs_reg_2_ ( .D(ns[2]), .CK(clk), .RN(rst_n), .Q(cs[2]) );
  DFFRHQX1 outset_cnt_reg_2_ ( .D(n5840), .CK(clk), .RN(rst_n), .Q(N944) );
  DFFRHQX1 calin_cnt_reg_0_ ( .D(N1362), .CK(clk), .RN(rst_n), .Q(calin_cnt[0]) );
  DFFRHQX1 store_cnt_reg_2_ ( .D(N14272), .CK(clk), .RN(rst_n), .Q(
        store_cnt[2]) );
  DFFRHQX1 cs_reg_1_ ( .D(ns[1]), .CK(clk), .RN(rst_n), .Q(cs[1]) );
  DFFRHQX1 cs_reg_0_ ( .D(ns[0]), .CK(clk), .RN(rst_n), .Q(cs[0]) );
  DFFRHQX1 m_size_reg_1_ ( .D(n4471), .CK(clk), .RN(rst_n), .Q(m_size[1]) );
  DFFRHQX1 out_value_reg ( .D(N14331), .CK(clk), .RN(rst_n), .Q(out_value) );
  DFFRHQX1 w_matrix_reg_1__0__15_ ( .D(n2540), .CK(clk), .RN(rst_n), .Q(
        w_matrix[895]) );
  DFFRHQX1 w_matrix_reg_1__0__13_ ( .D(n2542), .CK(clk), .RN(rst_n), .Q(
        w_matrix[893]) );
  DFFRHQX1 w_matrix_reg_1__0__12_ ( .D(n2543), .CK(clk), .RN(rst_n), .Q(
        w_matrix[892]) );
  DFFRHQX1 w_matrix_reg_1__0__11_ ( .D(n2544), .CK(clk), .RN(rst_n), .Q(
        w_matrix[891]) );
  DFFRHQX1 w_matrix_reg_1__0__10_ ( .D(n2545), .CK(clk), .RN(rst_n), .Q(
        w_matrix[890]) );
  DFFRHQX1 w_matrix_reg_1__0__9_ ( .D(n2546), .CK(clk), .RN(rst_n), .Q(
        w_matrix[889]) );
  DFFRHQX1 w_matrix_reg_1__0__8_ ( .D(n2547), .CK(clk), .RN(rst_n), .Q(
        w_matrix[888]) );
  DFFRHQX1 w_matrix_reg_1__0__7_ ( .D(n2548), .CK(clk), .RN(rst_n), .Q(
        w_matrix[887]) );
  DFFRHQX1 w_matrix_reg_1__0__6_ ( .D(n2549), .CK(clk), .RN(rst_n), .Q(
        w_matrix[886]) );
  DFFRHQX1 w_matrix_reg_1__0__5_ ( .D(n2550), .CK(clk), .RN(rst_n), .Q(
        w_matrix[885]) );
  DFFRHQX1 w_matrix_reg_1__0__4_ ( .D(n2551), .CK(clk), .RN(rst_n), .Q(
        w_matrix[884]) );
  DFFRHQX1 w_matrix_reg_1__0__3_ ( .D(n2552), .CK(clk), .RN(rst_n), .Q(
        w_matrix[883]) );
  DFFRHQX1 w_matrix_reg_1__0__2_ ( .D(n2553), .CK(clk), .RN(rst_n), .Q(
        w_matrix[882]) );
  DFFRHQX1 w_matrix_reg_1__0__1_ ( .D(n2554), .CK(clk), .RN(rst_n), .Q(
        w_matrix[881]) );
  DFFRHQX1 calweight_addr_reg_5_ ( .D(n5817), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[5]) );
  DFFRHQX1 calweight_addr_reg_6_ ( .D(n5818), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[6]) );
  DFFRHQX1 calweight_addr_reg_7_ ( .D(n5819), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[7]) );
  DFFRHQX1 calin_addr_reg_5_ ( .D(n5808), .CK(clk), .RN(rst_n), .Q(
        calin_addr[5]) );
  DFFRHQX1 calin_addr_reg_6_ ( .D(n5809), .CK(clk), .RN(rst_n), .Q(
        calin_addr[6]) );
  DFFRHQX1 calin_addr_reg_7_ ( .D(n5810), .CK(clk), .RN(rst_n), .Q(
        calin_addr[7]) );
  DFFRHQX1 cal_cnt_reg_4_ ( .D(N11318), .CK(clk), .RN(rst_n), .Q(cal_cnt[4])
         );
  DFFRHQX1 calweight_addr_reg_1_ ( .D(n5813), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[1]) );
  DFFRHQX1 calweight_addr_reg_2_ ( .D(n5814), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[2]) );
  DFFRHQX1 calweight_addr_reg_3_ ( .D(n5815), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[3]) );
  DFFRHQX1 calweight_addr_reg_4_ ( .D(n5816), .CK(clk), .RN(rst_n), .Q(
        calweight_addr[4]) );
  DFFRHQX1 calin_addr_reg_1_ ( .D(n5804), .CK(clk), .RN(rst_n), .Q(
        calin_addr[1]) );
  DFFRHQX1 calin_addr_reg_2_ ( .D(n5805), .CK(clk), .RN(rst_n), .Q(
        calin_addr[2]) );
  DFFRHQX1 calin_addr_reg_3_ ( .D(n5806), .CK(clk), .RN(rst_n), .Q(
        calin_addr[3]) );
  DFFRHQX1 calin_addr_reg_4_ ( .D(n5807), .CK(clk), .RN(rst_n), .Q(
        calin_addr[4]) );
  DFFRHQX1 c_plus_reg_5_ ( .D(N12571), .CK(clk), .RN(rst_n), .Q(c_plus[5]) );
  DFFRHQX1 c_plus_reg_4_ ( .D(N12570), .CK(clk), .RN(rst_n), .Q(c_plus[4]) );
  DFFRHQX1 cal_cnt_reg_5_ ( .D(N11319), .CK(clk), .RN(rst_n), .Q(cal_cnt[5])
         );
  DFFRHQX1 cal_cnt_reg_6_ ( .D(N11320), .CK(clk), .RN(rst_n), .Q(cal_cnt[6])
         );
  DFFRHQX1 c_plus_reg_13_ ( .D(N12579), .CK(clk), .RN(rst_n), .Q(c_plus[13])
         );
  DFFRHQX1 calin_cnt_reg_6_ ( .D(N1368), .CK(clk), .RN(rst_n), .Q(calin_cnt[6]) );
  DFFRHQX1 calin_cnt_reg_5_ ( .D(N1367), .CK(clk), .RN(rst_n), .Q(calin_cnt[5]) );
  DFFRHQX1 calin_cnt_reg_4_ ( .D(N1366), .CK(clk), .RN(rst_n), .Q(calin_cnt[4]) );
  JKFFRXL outset_cnt_reg_1_ ( .J(n741), .K(n743), .CK(clk), .RN(rst_n), .Q(
        N943), .QN(n4489) );
  DFFRHQX1 cs_reg_3_ ( .D(n5841), .CK(clk), .RN(rst_n), .Q(cs[3]) );
  DFFRHQX1 c_plus_reg_27_ ( .D(N12593), .CK(clk), .RN(rst_n), .Q(c_plus[27])
         );
  DFFRHQX1 c_plus_reg_22_ ( .D(N12588), .CK(clk), .RN(rst_n), .Q(c_plus[22])
         );
  DFFRHQX1 c_plus_reg_28_ ( .D(N12594), .CK(clk), .RN(rst_n), .Q(c_plus[28])
         );
  DFFRHQX1 c_plus_reg_16_ ( .D(N12582), .CK(clk), .RN(rst_n), .Q(c_plus[16])
         );
  DFFRHQX1 c_plus_reg_20_ ( .D(N12586), .CK(clk), .RN(rst_n), .Q(c_plus[20])
         );
  DFFRHQX1 c_plus_reg_15_ ( .D(N12581), .CK(clk), .RN(rst_n), .Q(c_plus[15])
         );
  DFFRHQX1 c_plus_reg_23_ ( .D(N12589), .CK(clk), .RN(rst_n), .Q(c_plus[23])
         );
  DFFRHQX1 store_cnt_reg_1_ ( .D(N14271), .CK(clk), .RN(rst_n), .Q(
        store_cnt[1]) );
  DFFRHQX1 calin_cnt_reg_3_ ( .D(N1365), .CK(clk), .RN(rst_n), .Q(calin_cnt[3]) );
  DFFRHQX1 c_plus_reg_37_ ( .D(N12603), .CK(clk), .RN(rst_n), .Q(c_plus[37])
         );
  DFFRHQX1 c_plus_reg_34_ ( .D(N12600), .CK(clk), .RN(rst_n), .Q(c_plus[34])
         );
  DFFRHQX1 c_plus_reg_38_ ( .D(N12604), .CK(clk), .RN(rst_n), .Q(c_plus[38])
         );
  DFFRHQX1 c_plus_reg_35_ ( .D(N12601), .CK(clk), .RN(rst_n), .Q(c_plus[35])
         );
  DFFRHQX1 out_valid_reg ( .D(n5878), .CK(clk), .RN(rst_n), .Q(out_valid) );
  DFFRHQX2 calin_cnt_reg_2_ ( .D(N1364), .CK(clk), .RN(rst_n), .Q(calin_cnt[2]) );
  DFFRHQX2 cal_cnt_reg_0_ ( .D(N11314), .CK(clk), .RN(rst_n), .Q(cal_cnt[0])
         );
  DFFRHQX1 out_cnt_reg_2_ ( .D(n5837), .CK(clk), .RN(rst_n), .Q(out_cnt[2]) );
  DFFRHQX1 store_cnt_reg_0_ ( .D(N14270), .CK(clk), .RN(rst_n), .Q(
        store_cnt[0]) );
  NOR2X1 U4358 ( .A(n873), .B(store_cnt[3]), .Y(n867) );
  AOI22X1 U4359 ( .A0(calin_cnt[2]), .A1(n5061), .B0(n5064), .B1(calin_cnt[3]), 
        .Y(n936) );
  AOI22X1 U4360 ( .A0(calin_cnt[1]), .A1(n5061), .B0(n5064), .B1(calin_cnt[2]), 
        .Y(n937) );
  AOI22X1 U4361 ( .A0(calin_cnt[0]), .A1(n5061), .B0(n5064), .B1(calin_cnt[1]), 
        .Y(n951) );
  AOI222XL U4362 ( .A0(value_out[25]), .A1(n1062), .B0(value_out[27]), .B1(
        n1060), .C0(value_out[26]), .C1(n1061), .Y(n1068) );
  NOR2X2 U4363 ( .A(n5971), .B(out_cnt[1]), .Y(n1062) );
  INVX1 U4364 ( .A(n882), .Y(n5895) );
  NAND2X1 U4365 ( .A(n867), .B(store_cnt[2]), .Y(n869) );
  NOR4X1 U4366 ( .A(cal_cnt[5]), .B(cal_cnt[4]), .C(cal_cnt[7]), .D(cal_cnt[6]), .Y(n1648) );
  AOI221X1 U4367 ( .A0(c_plus[5]), .A1(n832), .B0(c_plus[37]), .B1(n5970), 
        .C0(n833), .Y(n831) );
  NOR2X1 U4368 ( .A(n923), .B(mem_num_0), .Y(n931) );
  NOR3X2 U4369 ( .A(n728), .B(N14321), .C(n726), .Y(n753) );
  NAND2BX1 U4370 ( .AN(store_cnt[0]), .B(store_cnt[1]), .Y(n864) );
  NAND2BX1 U4371 ( .AN(store_cnt[1]), .B(store_cnt[0]), .Y(n862) );
  AOI22X2 U4372 ( .A0(n1038), .A1(n5050), .B0(n5878), .B1(n1039), .Y(n754) );
  NOR3X1 U4373 ( .A(n728), .B(n727), .C(n726), .Y(n1012) );
  AOI222X1 U4374 ( .A0(length_out[2]), .A1(N14321), .B0(n1088), .B1(
        length_out[0]), .C0(length_out[4]), .C1(n1089), .Y(n1086) );
  AOI222X1 U4375 ( .A0(length_out[3]), .A1(N14321), .B0(n1088), .B1(
        length_out[1]), .C0(length_out[5]), .C1(n1089), .Y(n1087) );
  INVX1 U4376 ( .A(cs[2]), .Y(n5889) );
  INVX1 U4377 ( .A(cs[3]), .Y(n5858) );
  NAND4X2 U4378 ( .A(cs[2]), .B(cs[0]), .C(n5890), .D(n5858), .Y(n873) );
  NAND4X2 U4379 ( .A(cs[3]), .B(n5883), .C(n5890), .D(n5889), .Y(n746) );
  NAND2X1 U4380 ( .A(store_cnt[1]), .B(store_cnt[0]), .Y(n866) );
  BUFX3 U4381 ( .A(n1516), .Y(n5056) );
  BUFX3 U4382 ( .A(n1450), .Y(n5055) );
  BUFX3 U4383 ( .A(n1583), .Y(n5053) );
  BUFX3 U4384 ( .A(n1651), .Y(n5054) );
  CLKINVX3 U4385 ( .A(c_plus[2]), .Y(n5932) );
  CLKINVX3 U4386 ( .A(c_plus[30]), .Y(n5962) );
  CLKINVX3 U4387 ( .A(c_plus[16]), .Y(n5947) );
  CLKINVX3 U4388 ( .A(c_plus[15]), .Y(n5946) );
  CLKINVX3 U4389 ( .A(c_plus[14]), .Y(n5945) );
  CLKINVX3 U4390 ( .A(c_plus[9]), .Y(n5939) );
  CLKINVX3 U4391 ( .A(c_plus[6]), .Y(n5936) );
  CLKINVX3 U4392 ( .A(c_plus[4]), .Y(n5934) );
  CLKINVX3 U4393 ( .A(c_plus[1]), .Y(n5931) );
  CLKINVX3 U4394 ( .A(c_plus[0]), .Y(n5930) );
  NAND4X2 U4395 ( .A(n1122), .B(n1121), .C(n1123), .D(n1124), .Y(ns[0]) );
  NAND4BXL U4396 ( .AN(calin_cnt[4]), .B(n1130), .C(n1131), .D(n1132), .Y(
        n1122) );
  NAND3BX2 U4397 ( .AN(n1115), .B(n1117), .C(n5066), .Y(ns[1]) );
  AOI22X1 U4398 ( .A0(n5053), .A1(x_matrix[641]), .B0(n5054), .B1(
        x_matrix[753]), .Y(n1710) );
  AOI22X1 U4399 ( .A0(n5055), .A1(x_matrix[433]), .B0(n5056), .B1(
        x_matrix[529]), .Y(n1711) );
  AOI22X1 U4400 ( .A0(n5053), .A1(x_matrix[643]), .B0(n5054), .B1(
        x_matrix[755]), .Y(n1702) );
  AOI22X1 U4401 ( .A0(n5055), .A1(x_matrix[435]), .B0(n5056), .B1(
        x_matrix[531]), .Y(n1703) );
  AOI22X1 U4402 ( .A0(n5053), .A1(x_matrix[640]), .B0(n5054), .B1(
        x_matrix[752]), .Y(n1714) );
  AOI22X1 U4403 ( .A0(n5055), .A1(x_matrix[432]), .B0(n5056), .B1(
        x_matrix[528]), .Y(n1715) );
  AOI22X1 U4404 ( .A0(n5053), .A1(x_matrix[645]), .B0(n5054), .B1(
        x_matrix[757]), .Y(n1694) );
  AOI22X1 U4405 ( .A0(n5055), .A1(x_matrix[437]), .B0(n5056), .B1(
        x_matrix[533]), .Y(n1695) );
  AOI22X1 U4406 ( .A0(n5053), .A1(x_matrix[647]), .B0(n5054), .B1(
        x_matrix[759]), .Y(n1686) );
  AOI22X1 U4407 ( .A0(n5055), .A1(x_matrix[439]), .B0(n5056), .B1(
        x_matrix[535]), .Y(n1687) );
  AOI22X1 U4408 ( .A0(n5053), .A1(x_matrix[649]), .B0(n5054), .B1(
        x_matrix[761]), .Y(n1678) );
  AOI22X1 U4409 ( .A0(n5055), .A1(x_matrix[441]), .B0(n5056), .B1(
        x_matrix[537]), .Y(n1679) );
  AOI22X1 U4410 ( .A0(n5053), .A1(x_matrix[642]), .B0(n5054), .B1(
        x_matrix[754]), .Y(n1706) );
  AOI22X1 U4411 ( .A0(n5055), .A1(x_matrix[434]), .B0(n5056), .B1(
        x_matrix[530]), .Y(n1707) );
  AOI22X1 U4412 ( .A0(n5053), .A1(x_matrix[644]), .B0(n5054), .B1(
        x_matrix[756]), .Y(n1698) );
  AOI22X1 U4413 ( .A0(n5055), .A1(x_matrix[436]), .B0(n5056), .B1(
        x_matrix[532]), .Y(n1699) );
  AOI22X1 U4414 ( .A0(n5053), .A1(x_matrix[646]), .B0(n5054), .B1(
        x_matrix[758]), .Y(n1690) );
  AOI22X1 U4415 ( .A0(n5055), .A1(x_matrix[438]), .B0(n5056), .B1(
        x_matrix[534]), .Y(n1691) );
  AOI22X1 U4416 ( .A0(n5053), .A1(x_matrix[651]), .B0(n5054), .B1(
        x_matrix[763]), .Y(n1670) );
  AOI22X1 U4417 ( .A0(n5055), .A1(x_matrix[443]), .B0(n5056), .B1(
        x_matrix[539]), .Y(n1671) );
  AOI31XL U4418 ( .A0(n1662), .A1(n1663), .A2(n1664), .B0(n1656), .Y(N11407)
         );
  AOI22X1 U4419 ( .A0(n5053), .A1(x_matrix[653]), .B0(n5054), .B1(
        x_matrix[765]), .Y(n1662) );
  AOI22X1 U4420 ( .A0(n5055), .A1(x_matrix[445]), .B0(n5056), .B1(
        x_matrix[541]), .Y(n1663) );
  AOI31X1 U4421 ( .A0(n1682), .A1(n1683), .A2(n1684), .B0(n1656), .Y(N11402)
         );
  AOI22X1 U4422 ( .A0(n5053), .A1(x_matrix[648]), .B0(n5054), .B1(
        x_matrix[760]), .Y(n1682) );
  AOI22X1 U4423 ( .A0(n5055), .A1(x_matrix[440]), .B0(n5056), .B1(
        x_matrix[536]), .Y(n1683) );
  AOI31X1 U4424 ( .A0(n1674), .A1(n1675), .A2(n1676), .B0(n1656), .Y(N11404)
         );
  AOI22X1 U4425 ( .A0(n5053), .A1(x_matrix[650]), .B0(n5054), .B1(
        x_matrix[762]), .Y(n1674) );
  AOI221XL U4426 ( .A0(n1318), .A1(x_matrix[250]), .B0(n1384), .B1(
        x_matrix[346]), .C0(n1677), .Y(n1676) );
  AOI22X1 U4427 ( .A0(n5055), .A1(x_matrix[442]), .B0(n5056), .B1(
        x_matrix[538]), .Y(n1675) );
  AOI31X1 U4428 ( .A0(n1666), .A1(n1667), .A2(n1668), .B0(n1656), .Y(N11406)
         );
  AOI22X1 U4429 ( .A0(n5053), .A1(x_matrix[652]), .B0(n5054), .B1(
        x_matrix[764]), .Y(n1666) );
  AOI221XL U4430 ( .A0(n1318), .A1(x_matrix[252]), .B0(n1384), .B1(
        x_matrix[348]), .C0(n1669), .Y(n1668) );
  AOI22X1 U4431 ( .A0(n5055), .A1(x_matrix[444]), .B0(n5056), .B1(
        x_matrix[540]), .Y(n1667) );
  AOI31X1 U4432 ( .A0(n1653), .A1(n1654), .A2(n1655), .B0(n1656), .Y(N11409)
         );
  AOI22X1 U4433 ( .A0(n5053), .A1(x_matrix[655]), .B0(n5054), .B1(
        x_matrix[767]), .Y(n1653) );
  AOI221X1 U4434 ( .A0(n1318), .A1(x_matrix[255]), .B0(n1384), .B1(
        x_matrix[351]), .C0(n1657), .Y(n1655) );
  AOI22X1 U4435 ( .A0(n5055), .A1(x_matrix[447]), .B0(n5056), .B1(
        x_matrix[543]), .Y(n1654) );
  AOI31X1 U4436 ( .A0(n1658), .A1(n1659), .A2(n1660), .B0(n1656), .Y(N11408)
         );
  AOI22X1 U4437 ( .A0(n5053), .A1(x_matrix[654]), .B0(n5054), .B1(
        x_matrix[766]), .Y(n1658) );
  AOI221X1 U4438 ( .A0(n1318), .A1(x_matrix[254]), .B0(n1384), .B1(
        x_matrix[350]), .C0(n1661), .Y(n1660) );
  AOI22X1 U4439 ( .A0(n5055), .A1(x_matrix[446]), .B0(n5056), .B1(
        x_matrix[542]), .Y(n1659) );
  NOR3X2 U4440 ( .A(ns[0]), .B(ns[1]), .C(n5823), .Y(n4473) );
  NOR3X2 U4441 ( .A(ns[0]), .B(ns[1]), .C(n5823), .Y(n4474) );
  OAI31X1 U4442 ( .A0(n939), .A1(n5859), .A2(n935), .B0(n925), .Y(n942) );
  OAI31X1 U4443 ( .A0(n939), .A1(n5859), .A2(n930), .B0(n925), .Y(n940) );
  OAI31X1 U4444 ( .A0(n939), .A1(n927), .A2(n5859), .B0(n925), .Y(n938) );
  AND2X2 U4445 ( .A(n4504), .B(n4508), .Y(n4881) );
  AND2X2 U4446 ( .A(n4499), .B(n4506), .Y(n4871) );
  AND2X2 U4447 ( .A(n4505), .B(n4508), .Y(n4880) );
  AND2X2 U4448 ( .A(n4498), .B(n4505), .Y(n4868) );
  AND2X2 U4449 ( .A(n4499), .B(n4505), .Y(n4872) );
  AND2X2 U4450 ( .A(n4507), .B(n4509), .Y(n4866) );
  AND2X2 U4451 ( .A(n4498), .B(n4509), .Y(n4870) );
  AND2X2 U4452 ( .A(n4507), .B(n4505), .Y(n4878) );
  AND2X2 U4453 ( .A(n4509), .B(n4508), .Y(n4883) );
  AND2X2 U4454 ( .A(mem_num_0), .B(n5050), .Y(n1138) );
  AND2X2 U4455 ( .A(n4499), .B(n4504), .Y(n4873) );
  AND2X2 U4456 ( .A(n4498), .B(n4506), .Y(n4867) );
  AND2X2 U4457 ( .A(n4498), .B(n4504), .Y(n4869) );
  AND2X2 U4458 ( .A(n4507), .B(n4504), .Y(n4879) );
  AND2X2 U4459 ( .A(n4507), .B(n4506), .Y(n4884) );
  INVX8 U4460 ( .A(n5315), .Y(n5314) );
  AND2X2 U4461 ( .A(n5050), .B(n884), .Y(n4475) );
  AND2X2 U4462 ( .A(n5050), .B(n883), .Y(n4476) );
  AND2X2 U4463 ( .A(n5050), .B(n880), .Y(n4477) );
  AND2X2 U4464 ( .A(n5050), .B(n878), .Y(n4478) );
  AND2X2 U4465 ( .A(n5050), .B(n877), .Y(n4479) );
  AND2X2 U4466 ( .A(n5050), .B(n876), .Y(n4480) );
  AND2X2 U4467 ( .A(n5050), .B(n874), .Y(n4481) );
  AND2X2 U4468 ( .A(n5050), .B(n872), .Y(n4482) );
  AND2X2 U4469 ( .A(n5050), .B(n871), .Y(n4483) );
  AND2X2 U4470 ( .A(n5050), .B(n870), .Y(n4484) );
  AND2X2 U4471 ( .A(n5050), .B(n868), .Y(n4485) );
  AND2X2 U4472 ( .A(n5050), .B(n865), .Y(n4486) );
  AND2X2 U4473 ( .A(n5050), .B(n863), .Y(n4487) );
  AND2X2 U4474 ( .A(n5050), .B(n861), .Y(n4488) );
  OAI31X1 U4475 ( .A0(n949), .A1(n5859), .A2(n935), .B0(n925), .Y(n957) );
  OAI31X1 U4476 ( .A0(n949), .A1(n5859), .A2(n930), .B0(n925), .Y(n952) );
  OAI31X1 U4477 ( .A0(n939), .A1(n5859), .A2(n933), .B0(n925), .Y(n941) );
  NAND3X2 U4478 ( .A(n1118), .B(n5890), .C(cs[2]), .Y(n923) );
  NOR2X1 U4479 ( .A(n5058), .B(n5086), .Y(n1254) );
  NOR2X2 U4480 ( .A(m_size[1]), .B(m_size[0]), .Y(mem_num_0) );
  CLKINVX3 U4481 ( .A(n923), .Y(n5249) );
  INVX1 U4482 ( .A(n5563), .Y(n5559) );
  INVX1 U4483 ( .A(n5380), .Y(n5379) );
  INVX1 U4484 ( .A(n5402), .Y(n5401) );
  NAND2X1 U4485 ( .A(n5249), .B(n5073), .Y(n917) );
  NAND2X1 U4486 ( .A(n5249), .B(n5074), .Y(n916) );
  NAND2X1 U4487 ( .A(n5249), .B(n5075), .Y(n915) );
  NAND2X1 U4488 ( .A(n5249), .B(n5076), .Y(n914) );
  NAND2X1 U4489 ( .A(n5249), .B(n5077), .Y(n909) );
  NAND2X1 U4490 ( .A(n5249), .B(n5078), .Y(n887) );
  NAND2X1 U4491 ( .A(n5249), .B(n941), .Y(n912) );
  NAND2X1 U4492 ( .A(n5249), .B(n938), .Y(n910) );
  NAND2X1 U4493 ( .A(n5250), .B(n957), .Y(n921) );
  NAND2X1 U4494 ( .A(n5250), .B(n952), .Y(n919) );
  NAND2X1 U4495 ( .A(n5250), .B(n5071), .Y(n920) );
  NAND2X1 U4496 ( .A(n5250), .B(n5072), .Y(n918) );
  NAND2X1 U4497 ( .A(n5249), .B(n5378), .Y(n913) );
  NAND2X1 U4498 ( .A(n5249), .B(n5400), .Y(n911) );
  INVX1 U4499 ( .A(n5071), .Y(n5337) );
  INVX1 U4500 ( .A(n5072), .Y(n5350) );
  INVX1 U4501 ( .A(n957), .Y(n5799) );
  INVX1 U4502 ( .A(n952), .Y(n5800) );
  INVX1 U4503 ( .A(n938), .Y(n5802) );
  INVX1 U4504 ( .A(n941), .Y(n5801) );
  AOI21X1 U4505 ( .A0(n931), .A1(n932), .B0(n5797), .Y(n908) );
  OAI21XL U4506 ( .A0(n924), .A1(n5859), .B0(n925), .Y(n926) );
  NAND3X1 U4507 ( .A(n5569), .B(n907), .C(n925), .Y(n906) );
  CLKINVX3 U4508 ( .A(n923), .Y(n5250) );
  NOR2X1 U4509 ( .A(n933), .B(n928), .Y(n932) );
  OAI21XL U4510 ( .A0(n5895), .A1(n875), .B0(n5065), .Y(n874) );
  OAI21XL U4511 ( .A0(n5895), .A1(n859), .B0(n5065), .Y(n858) );
  INVX1 U4512 ( .A(ns[0]), .Y(n5821) );
  INVX1 U4513 ( .A(ns[1]), .Y(n5822) );
  NOR2X1 U4514 ( .A(n5061), .B(n5064), .Y(n1128) );
  BUFX3 U4515 ( .A(n5842), .Y(n5050) );
  NAND2X1 U4516 ( .A(n5053), .B(n5086), .Y(n1257) );
  NAND4X1 U4517 ( .A(n1044), .B(n5975), .C(n5976), .D(n5977), .Y(n755) );
  NAND2X1 U4518 ( .A(n1648), .B(n1649), .Y(n1182) );
  INVX1 U4519 ( .A(n746), .Y(n5878) );
  INVX1 U4520 ( .A(n951), .Y(n5880) );
  NAND2X1 U4521 ( .A(n867), .B(n5896), .Y(n859) );
  NAND2X1 U4522 ( .A(n879), .B(n5896), .Y(n875) );
  NAND2X1 U4523 ( .A(n5054), .B(n5086), .Y(n1185) );
  NOR2X1 U4524 ( .A(n873), .B(n5897), .Y(n879) );
  OAI21XL U4525 ( .A0(n866), .A1(n875), .B0(n5065), .Y(n878) );
  OAI21XL U4526 ( .A0(n866), .A1(n869), .B0(n5065), .Y(n872) );
  OAI21XL U4527 ( .A0(n859), .A1(n866), .B0(n5065), .Y(n865) );
  OAI21XL U4528 ( .A0(n864), .A1(n881), .B0(n5065), .Y(n884) );
  OAI21XL U4529 ( .A0(n864), .A1(n875), .B0(n5065), .Y(n877) );
  OAI21XL U4530 ( .A0(n864), .A1(n869), .B0(n5065), .Y(n871) );
  OAI21XL U4531 ( .A0(n862), .A1(n881), .B0(n5065), .Y(n883) );
  OAI21XL U4532 ( .A0(n5895), .A1(n881), .B0(n5065), .Y(n880) );
  OAI21XL U4533 ( .A0(n859), .A1(n864), .B0(n5065), .Y(n863) );
  OAI21XL U4534 ( .A0(n859), .A1(n862), .B0(n5065), .Y(n861) );
  OAI21XL U4535 ( .A0(n862), .A1(n875), .B0(n5065), .Y(n876) );
  OAI21XL U4536 ( .A0(n862), .A1(n869), .B0(n5065), .Y(n870) );
  OAI21XL U4537 ( .A0(n5895), .A1(n869), .B0(n5065), .Y(n868) );
  INVX1 U4538 ( .A(n5086), .Y(n5894) );
  INVX1 U4539 ( .A(n5066), .Y(n5877) );
  OAI21XL U4540 ( .A0(n1009), .A1(n1010), .B0(in_valid), .Y(n1002) );
  CLKINVX3 U4541 ( .A(c_plus[33]), .Y(n5964) );
  CLKINVX3 U4542 ( .A(c_plus[32]), .Y(n5963) );
  CLKINVX3 U4543 ( .A(c_plus[36]), .Y(n5967) );
  NOR3X1 U4544 ( .A(c_plus[38]), .B(c_plus[39]), .C(c_plus[37]), .Y(n779) );
  NAND4X1 U4545 ( .A(n791), .B(n782), .C(n806), .D(n852), .Y(n826) );
  NAND4X1 U4546 ( .A(cs[0]), .B(cs[1]), .C(n5889), .D(n5858), .Y(n1121) );
  INVX1 U4547 ( .A(store_cnt[2]), .Y(n5896) );
  CLKINVX3 U4548 ( .A(c_plus[25]), .Y(n5957) );
  CLKINVX3 U4549 ( .A(c_plus[26]), .Y(n5958) );
  CLKINVX3 U4550 ( .A(c_plus[24]), .Y(n5955) );
  NOR2X1 U4551 ( .A(store_cnt[0]), .B(store_cnt[1]), .Y(n882) );
  CLKINVX3 U4552 ( .A(c_plus[29]), .Y(n5961) );
  NOR3X1 U4553 ( .A(c_plus[16]), .B(c_plus[17]), .C(c_plus[15]), .Y(n851) );
  NOR3X1 U4554 ( .A(n1043), .B(n755), .C(n5973), .Y(n1042) );
  NAND2X1 U4555 ( .A(c_plus[9]), .B(n829), .Y(n799) );
  NAND3X1 U4556 ( .A(n829), .B(n5939), .C(c_plus[8]), .Y(n801) );
  NAND3X1 U4557 ( .A(n834), .B(n835), .C(c_plus[13]), .Y(n816) );
  INVX1 U4558 ( .A(cs[0]), .Y(n5883) );
  BUFX3 U4559 ( .A(n5790), .Y(n5048) );
  BUFX3 U4560 ( .A(n5789), .Y(n5047) );
  BUFX3 U4561 ( .A(n5788), .Y(n5046) );
  BUFX3 U4562 ( .A(n5787), .Y(n5045) );
  BUFX3 U4563 ( .A(n5786), .Y(n5044) );
  BUFX3 U4564 ( .A(n5785), .Y(n5043) );
  BUFX3 U4565 ( .A(n5780), .Y(n5038) );
  BUFX3 U4566 ( .A(n5769), .Y(n5027) );
  BUFX3 U4567 ( .A(n5758), .Y(n5016) );
  BUFX3 U4568 ( .A(n5747), .Y(n5005) );
  BUFX3 U4569 ( .A(n5736), .Y(n4994) );
  BUFX3 U4570 ( .A(n5731), .Y(n4989) );
  BUFX3 U4571 ( .A(n5730), .Y(n4988) );
  BUFX3 U4572 ( .A(n5729), .Y(n4987) );
  BUFX3 U4573 ( .A(n5728), .Y(n4986) );
  CLKINVX3 U4574 ( .A(c_plus[21]), .Y(n5952) );
  CLKINVX3 U4575 ( .A(c_plus[11]), .Y(n5942) );
  BUFX3 U4576 ( .A(n5784), .Y(n5042) );
  BUFX3 U4577 ( .A(n5783), .Y(n5041) );
  BUFX3 U4578 ( .A(n5782), .Y(n5040) );
  BUFX3 U4579 ( .A(n5781), .Y(n5039) );
  BUFX3 U4580 ( .A(n5779), .Y(n5037) );
  BUFX3 U4581 ( .A(n5778), .Y(n5036) );
  BUFX3 U4582 ( .A(n5777), .Y(n5035) );
  BUFX3 U4583 ( .A(n5776), .Y(n5034) );
  BUFX3 U4584 ( .A(n5775), .Y(n5033) );
  BUFX3 U4585 ( .A(n5774), .Y(n5032) );
  BUFX3 U4586 ( .A(n5773), .Y(n5031) );
  BUFX3 U4587 ( .A(n5772), .Y(n5030) );
  BUFX3 U4588 ( .A(n5771), .Y(n5029) );
  BUFX3 U4589 ( .A(n5770), .Y(n5028) );
  BUFX3 U4590 ( .A(n5768), .Y(n5026) );
  BUFX3 U4591 ( .A(n5767), .Y(n5025) );
  BUFX3 U4592 ( .A(n5791), .Y(n5049) );
  CLKINVX3 U4593 ( .A(c_plus[8]), .Y(n5938) );
  CLKINVX3 U4594 ( .A(c_plus[10]), .Y(n5940) );
  CLKINVX3 U4595 ( .A(c_plus[12]), .Y(n5943) );
  BUFX3 U4596 ( .A(n5765), .Y(n5023) );
  BUFX3 U4597 ( .A(n5764), .Y(n5022) );
  BUFX3 U4598 ( .A(n5763), .Y(n5021) );
  BUFX3 U4599 ( .A(n5762), .Y(n5020) );
  BUFX3 U4600 ( .A(n5761), .Y(n5019) );
  BUFX3 U4601 ( .A(n5760), .Y(n5018) );
  BUFX3 U4602 ( .A(n5759), .Y(n5017) );
  BUFX3 U4603 ( .A(n5757), .Y(n5015) );
  BUFX3 U4604 ( .A(n5756), .Y(n5014) );
  BUFX3 U4605 ( .A(n5755), .Y(n5013) );
  BUFX3 U4606 ( .A(n5754), .Y(n5012) );
  BUFX3 U4607 ( .A(n5753), .Y(n5011) );
  BUFX3 U4608 ( .A(n5752), .Y(n5010) );
  BUFX3 U4609 ( .A(n5751), .Y(n5009) );
  BUFX3 U4610 ( .A(n5750), .Y(n5008) );
  BUFX3 U4611 ( .A(n5766), .Y(n5024) );
  BUFX3 U4612 ( .A(n5749), .Y(n5007) );
  BUFX3 U4613 ( .A(n5748), .Y(n5006) );
  BUFX3 U4614 ( .A(n5746), .Y(n5004) );
  BUFX3 U4615 ( .A(n5745), .Y(n5003) );
  BUFX3 U4616 ( .A(n5744), .Y(n5002) );
  BUFX3 U4617 ( .A(n5743), .Y(n5001) );
  BUFX3 U4618 ( .A(n5742), .Y(n5000) );
  BUFX3 U4619 ( .A(n5741), .Y(n4999) );
  BUFX3 U4620 ( .A(n5740), .Y(n4998) );
  BUFX3 U4621 ( .A(n5739), .Y(n4997) );
  BUFX3 U4622 ( .A(n5738), .Y(n4996) );
  BUFX3 U4623 ( .A(n5737), .Y(n4995) );
  BUFX3 U4624 ( .A(n5735), .Y(n4993) );
  BUFX3 U4625 ( .A(n5734), .Y(n4992) );
  BUFX3 U4626 ( .A(n5733), .Y(n4991) );
  BUFX3 U4627 ( .A(n5732), .Y(n4990) );
  BUFX3 U4628 ( .A(n5727), .Y(n4985) );
  BUFX3 U4629 ( .A(n5726), .Y(n4984) );
  BUFX3 U4630 ( .A(n5725), .Y(n4983) );
  BUFX3 U4631 ( .A(n5724), .Y(n4982) );
  BUFX3 U4632 ( .A(n5723), .Y(n4981) );
  BUFX3 U4633 ( .A(n5722), .Y(n4980) );
  BUFX3 U4634 ( .A(n5721), .Y(n4979) );
  BUFX3 U4635 ( .A(n5716), .Y(n4974) );
  BUFX3 U4636 ( .A(n5705), .Y(n4963) );
  BUFX3 U4637 ( .A(n5694), .Y(n4952) );
  BUFX3 U4638 ( .A(n5683), .Y(n4941) );
  BUFX3 U4639 ( .A(n5672), .Y(n4930) );
  BUFX3 U4640 ( .A(n5667), .Y(n4925) );
  BUFX3 U4641 ( .A(n5666), .Y(n4924) );
  BUFX3 U4642 ( .A(n5665), .Y(n4923) );
  BUFX3 U4643 ( .A(n5664), .Y(n4922) );
  BUFX3 U4644 ( .A(n5720), .Y(n4978) );
  BUFX3 U4645 ( .A(n5719), .Y(n4977) );
  BUFX3 U4646 ( .A(n5718), .Y(n4976) );
  BUFX3 U4647 ( .A(n5717), .Y(n4975) );
  BUFX3 U4648 ( .A(n5715), .Y(n4973) );
  BUFX3 U4649 ( .A(n5714), .Y(n4972) );
  BUFX3 U4650 ( .A(n5713), .Y(n4971) );
  BUFX3 U4651 ( .A(n5712), .Y(n4970) );
  BUFX3 U4652 ( .A(n5711), .Y(n4969) );
  BUFX3 U4653 ( .A(n5710), .Y(n4968) );
  BUFX3 U4654 ( .A(n5709), .Y(n4967) );
  BUFX3 U4655 ( .A(n5708), .Y(n4966) );
  BUFX3 U4656 ( .A(n5707), .Y(n4965) );
  BUFX3 U4657 ( .A(n5706), .Y(n4964) );
  BUFX3 U4658 ( .A(n5704), .Y(n4962) );
  BUFX3 U4659 ( .A(n5703), .Y(n4961) );
  BUFX3 U4660 ( .A(n5685), .Y(n4943) );
  BUFX3 U4661 ( .A(n5684), .Y(n4942) );
  BUFX3 U4662 ( .A(n5682), .Y(n4940) );
  BUFX3 U4663 ( .A(n5681), .Y(n4939) );
  BUFX3 U4664 ( .A(n5680), .Y(n4938) );
  BUFX3 U4665 ( .A(n5679), .Y(n4937) );
  BUFX3 U4666 ( .A(n5678), .Y(n4936) );
  BUFX3 U4667 ( .A(n5677), .Y(n4935) );
  BUFX3 U4668 ( .A(n5676), .Y(n4934) );
  BUFX3 U4669 ( .A(n5675), .Y(n4933) );
  BUFX3 U4670 ( .A(n5674), .Y(n4932) );
  BUFX3 U4671 ( .A(n5673), .Y(n4931) );
  BUFX3 U4672 ( .A(n5671), .Y(n4929) );
  BUFX3 U4673 ( .A(n5670), .Y(n4928) );
  BUFX3 U4674 ( .A(n5669), .Y(n4927) );
  BUFX3 U4675 ( .A(n5668), .Y(n4926) );
  BUFX3 U4676 ( .A(n5702), .Y(n4960) );
  BUFX3 U4677 ( .A(n5701), .Y(n4959) );
  BUFX3 U4678 ( .A(n5700), .Y(n4958) );
  BUFX3 U4679 ( .A(n5699), .Y(n4957) );
  BUFX3 U4680 ( .A(n5698), .Y(n4956) );
  BUFX3 U4681 ( .A(n5697), .Y(n4955) );
  BUFX3 U4682 ( .A(n5696), .Y(n4954) );
  BUFX3 U4683 ( .A(n5695), .Y(n4953) );
  BUFX3 U4684 ( .A(n5693), .Y(n4951) );
  BUFX3 U4685 ( .A(n5692), .Y(n4950) );
  BUFX3 U4686 ( .A(n5691), .Y(n4949) );
  BUFX3 U4687 ( .A(n5690), .Y(n4948) );
  BUFX3 U4688 ( .A(n5689), .Y(n4947) );
  BUFX3 U4689 ( .A(n5688), .Y(n4946) );
  BUFX3 U4690 ( .A(n5687), .Y(n4945) );
  BUFX3 U4691 ( .A(n5686), .Y(n4944) );
  INVX1 U4692 ( .A(store_cnt[3]), .Y(n5897) );
  NAND2X1 U4693 ( .A(N14263), .B(n5050), .Y(n1092) );
  NOR3X1 U4694 ( .A(calin_cnt[5]), .B(calin_cnt[7]), .C(calin_cnt[6]), .Y(
        n1131) );
  INVX1 U4695 ( .A(cal_cnt[0]), .Y(n5891) );
  INVX1 U4696 ( .A(out_cnt[3]), .Y(n5975) );
  NAND4X1 U4697 ( .A(n1003), .B(n1004), .C(n1005), .D(n1006), .Y(n967) );
  NAND2X1 U4698 ( .A(c_plus[26]), .B(n830), .Y(n806) );
  INVX1 U4699 ( .A(out_cnt[4]), .Y(n5976) );
  NAND2X1 U4700 ( .A(c_plus[25]), .B(n830), .Y(n805) );
  INVX1 U4701 ( .A(out_cnt[5]), .Y(n5977) );
  INVX1 U4702 ( .A(out_cnt[2]), .Y(n5974) );
  NOR4BX1 U4703 ( .AN(n1517), .B(in_cnt_64[1]), .C(in_cnt_64[2]), .D(
        in_cnt_64[0]), .Y(n739) );
  CLKINVX3 U4704 ( .A(c_plus[17]), .Y(n5948) );
  NAND2X1 U4705 ( .A(n879), .B(store_cnt[2]), .Y(n881) );
  ADDHXL U4706 ( .A(in_matrix_cnt[3]), .B(add_250_carry[3]), .CO(
        add_250_carry[4]), .S(N1088) );
  CLKINVX3 U4707 ( .A(c_plus[3]), .Y(n5933) );
  CLKINVX3 U4708 ( .A(c_plus[37]), .Y(n5968) );
  CLKINVX3 U4709 ( .A(c_plus[38]), .Y(n5969) );
  CLKINVX3 U4710 ( .A(n5502), .Y(n5493) );
  CLKINVX3 U4711 ( .A(n5524), .Y(n5515) );
  CLKINVX3 U4712 ( .A(n5458), .Y(n5455) );
  CLKINVX3 U4713 ( .A(n5480), .Y(n5477) );
  CLKINVX3 U4714 ( .A(n5469), .Y(n5466) );
  CLKINVX3 U4715 ( .A(n5491), .Y(n5488) );
  CLKINVX3 U4716 ( .A(n5546), .Y(n5543) );
  CLKINVX3 U4717 ( .A(n5581), .Y(n5578) );
  CLKINVX3 U4718 ( .A(n5500), .Y(n5499) );
  CLKINVX3 U4719 ( .A(n5522), .Y(n5521) );
  CLKINVX3 U4720 ( .A(n5500), .Y(n5498) );
  CLKINVX3 U4721 ( .A(n5522), .Y(n5520) );
  CLKINVX3 U4722 ( .A(n5425), .Y(n5422) );
  CLKINVX3 U4723 ( .A(n5447), .Y(n5444) );
  CLKINVX3 U4724 ( .A(n5424), .Y(n5421) );
  CLKINVX3 U4725 ( .A(n5446), .Y(n5443) );
  CLKINVX3 U4726 ( .A(n5412), .Y(n5407) );
  CLKINVX3 U4727 ( .A(n5434), .Y(n5429) );
  CLKINVX3 U4728 ( .A(n5511), .Y(n5506) );
  CLKINVX3 U4729 ( .A(n5533), .Y(n5529) );
  CLKINVX3 U4730 ( .A(n5425), .Y(n5416) );
  CLKINVX3 U4731 ( .A(n5447), .Y(n5438) );
  CLKINVX3 U4732 ( .A(n5423), .Y(n5420) );
  CLKINVX3 U4733 ( .A(n5445), .Y(n5442) );
  CLKINVX3 U4734 ( .A(n5500), .Y(n5497) );
  CLKINVX3 U4735 ( .A(n5522), .Y(n5519) );
  CLKINVX3 U4736 ( .A(n5469), .Y(n5465) );
  CLKINVX3 U4737 ( .A(n5491), .Y(n5487) );
  CLKINVX3 U4738 ( .A(n5546), .Y(n5542) );
  CLKINVX3 U4739 ( .A(n5581), .Y(n5577) );
  CLKINVX3 U4740 ( .A(n5457), .Y(n5454) );
  CLKINVX3 U4741 ( .A(n5479), .Y(n5476) );
  CLKINVX3 U4742 ( .A(n5412), .Y(n5409) );
  CLKINVX3 U4743 ( .A(n5434), .Y(n5431) );
  CLKINVX3 U4744 ( .A(n5511), .Y(n5508) );
  CLKINVX3 U4745 ( .A(n5534), .Y(n5530) );
  CLKINVX3 U4746 ( .A(n5456), .Y(n5452) );
  CLKINVX3 U4747 ( .A(n5478), .Y(n5474) );
  CLKINVX3 U4748 ( .A(n5412), .Y(n5410) );
  CLKINVX3 U4749 ( .A(n5434), .Y(n5432) );
  CLKINVX3 U4750 ( .A(n5511), .Y(n5509) );
  CLKINVX3 U4751 ( .A(n5533), .Y(n5531) );
  CLKINVX3 U4752 ( .A(n5456), .Y(n5451) );
  CLKINVX3 U4753 ( .A(n5478), .Y(n5473) );
  CLKINVX3 U4754 ( .A(n5467), .Y(n5464) );
  CLKINVX3 U4755 ( .A(n5489), .Y(n5486) );
  CLKINVX3 U4756 ( .A(n5544), .Y(n5541) );
  CLKINVX3 U4757 ( .A(n5579), .Y(n5576) );
  CLKINVX3 U4758 ( .A(n5467), .Y(n5463) );
  CLKINVX3 U4759 ( .A(n5489), .Y(n5485) );
  CLKINVX3 U4760 ( .A(n5544), .Y(n5540) );
  CLKINVX3 U4761 ( .A(n5579), .Y(n5575) );
  CLKINVX3 U4762 ( .A(n5414), .Y(n5411) );
  CLKINVX3 U4763 ( .A(n5436), .Y(n5433) );
  CLKINVX3 U4764 ( .A(n5513), .Y(n5510) );
  CLKINVX3 U4765 ( .A(n5535), .Y(n5532) );
  CLKINVX3 U4766 ( .A(n5457), .Y(n5450) );
  CLKINVX3 U4767 ( .A(n5479), .Y(n5472) );
  CLKINVX3 U4768 ( .A(n5456), .Y(n5453) );
  CLKINVX3 U4769 ( .A(n5478), .Y(n5475) );
  CLKINVX3 U4770 ( .A(n5467), .Y(n5462) );
  CLKINVX3 U4771 ( .A(n5489), .Y(n5484) );
  CLKINVX3 U4772 ( .A(n5544), .Y(n5539) );
  CLKINVX3 U4773 ( .A(n5579), .Y(n5574) );
  CLKINVX3 U4774 ( .A(n5414), .Y(n5408) );
  CLKINVX3 U4775 ( .A(n5436), .Y(n5430) );
  CLKINVX3 U4776 ( .A(n5468), .Y(n5461) );
  CLKINVX3 U4777 ( .A(n5490), .Y(n5483) );
  CLKINVX3 U4778 ( .A(n5513), .Y(n5507) );
  CLKINVX3 U4779 ( .A(n5545), .Y(n5538) );
  CLKINVX3 U4780 ( .A(n5580), .Y(n5573) );
  CLKINVX3 U4781 ( .A(n5423), .Y(n5418) );
  CLKINVX3 U4782 ( .A(n5445), .Y(n5440) );
  CLKINVX3 U4783 ( .A(n5501), .Y(n5496) );
  CLKINVX3 U4784 ( .A(n5523), .Y(n5518) );
  CLKINVX3 U4785 ( .A(n5424), .Y(n5417) );
  CLKINVX3 U4786 ( .A(n5446), .Y(n5439) );
  CLKINVX3 U4787 ( .A(n5501), .Y(n5495) );
  CLKINVX3 U4788 ( .A(n5523), .Y(n5517) );
  CLKINVX3 U4789 ( .A(n5502), .Y(n5494) );
  CLKINVX3 U4790 ( .A(n5524), .Y(n5516) );
  CLKINVX3 U4791 ( .A(n5423), .Y(n5419) );
  CLKINVX3 U4792 ( .A(n5445), .Y(n5441) );
  CLKINVX3 U4793 ( .A(n5414), .Y(n5404) );
  CLKINVX3 U4794 ( .A(n5436), .Y(n5426) );
  CLKINVX3 U4795 ( .A(n5458), .Y(n5449) );
  CLKINVX3 U4796 ( .A(n5480), .Y(n5471) );
  CLKINVX3 U4797 ( .A(n5513), .Y(n5503) );
  CLKINVX3 U4798 ( .A(n5535), .Y(n5525) );
  CLKINVX3 U4799 ( .A(n5468), .Y(n5460) );
  CLKINVX3 U4800 ( .A(n5490), .Y(n5482) );
  CLKINVX3 U4801 ( .A(n5545), .Y(n5537) );
  CLKINVX3 U4802 ( .A(n5580), .Y(n5572) );
  CLKINVX3 U4803 ( .A(n5535), .Y(n5526) );
  CLKINVX3 U4804 ( .A(n5469), .Y(n5459) );
  CLKINVX3 U4805 ( .A(n5491), .Y(n5481) );
  CLKINVX3 U4806 ( .A(n5546), .Y(n5536) );
  CLKINVX3 U4807 ( .A(n5581), .Y(n5571) );
  CLKINVX3 U4808 ( .A(n5413), .Y(n5405) );
  CLKINVX3 U4809 ( .A(n5435), .Y(n5427) );
  CLKINVX3 U4810 ( .A(n5512), .Y(n5504) );
  CLKINVX3 U4811 ( .A(n5534), .Y(n5527) );
  CLKINVX3 U4812 ( .A(n5413), .Y(n5406) );
  CLKINVX3 U4813 ( .A(n5435), .Y(n5428) );
  CLKINVX3 U4814 ( .A(n5512), .Y(n5505) );
  CLKINVX3 U4815 ( .A(n5534), .Y(n5528) );
  CLKINVX3 U4816 ( .A(n5425), .Y(n5415) );
  CLKINVX3 U4817 ( .A(n5447), .Y(n5437) );
  CLKINVX3 U4818 ( .A(n5502), .Y(n5492) );
  CLKINVX3 U4819 ( .A(n5524), .Y(n5514) );
  CLKINVX3 U4820 ( .A(n5561), .Y(n5558) );
  INVX1 U4821 ( .A(n5379), .Y(n5362) );
  INVX1 U4822 ( .A(n5401), .Y(n5384) );
  INVX1 U4823 ( .A(n957), .Y(n5092) );
  INVX1 U4824 ( .A(n952), .Y(n5102) );
  INVX1 U4825 ( .A(n941), .Y(n5144) );
  INVX1 U4826 ( .A(n5160), .Y(n5155) );
  INVX1 U4827 ( .A(n5098), .Y(n5089) );
  INVX1 U4828 ( .A(n5108), .Y(n5099) );
  INVX1 U4829 ( .A(n5073), .Y(n5110) );
  INVX1 U4830 ( .A(n5075), .Y(n5126) );
  INVX1 U4831 ( .A(n5150), .Y(n5141) );
  INVX1 U4832 ( .A(n5160), .Y(n5152) );
  INVX1 U4833 ( .A(n5098), .Y(n5090) );
  INVX1 U4834 ( .A(n5108), .Y(n5100) );
  INVX1 U4835 ( .A(n947), .Y(n5111) );
  INVX1 U4836 ( .A(n945), .Y(n5127) );
  INVX1 U4837 ( .A(n5150), .Y(n5142) );
  INVX1 U4838 ( .A(n5160), .Y(n5153) );
  INVX1 U4839 ( .A(n5074), .Y(n5118) );
  INVX1 U4840 ( .A(n5076), .Y(n5133) );
  INVX1 U4841 ( .A(n5077), .Y(n5162) );
  INVX1 U4842 ( .A(n5078), .Y(n5170) );
  INVX1 U4843 ( .A(n5098), .Y(n5091) );
  INVX1 U4844 ( .A(n5108), .Y(n5101) );
  INVX1 U4845 ( .A(n5150), .Y(n5143) );
  INVX1 U4846 ( .A(n5076), .Y(n5134) );
  INVX1 U4847 ( .A(n5160), .Y(n5154) );
  INVX1 U4848 ( .A(n946), .Y(n5119) );
  INVX1 U4849 ( .A(n5076), .Y(n5135) );
  INVX1 U4850 ( .A(n934), .Y(n5163) );
  INVX1 U4851 ( .A(n929), .Y(n5171) );
  INVX1 U4852 ( .A(n5378), .Y(n5361) );
  INVX1 U4853 ( .A(n5400), .Y(n5383) );
  INVX1 U4854 ( .A(n5378), .Y(n5360) );
  INVX1 U4855 ( .A(n5400), .Y(n5382) );
  INVX1 U4856 ( .A(n5371), .Y(n5366) );
  INVX1 U4857 ( .A(n5393), .Y(n5388) );
  INVX1 U4858 ( .A(n5073), .Y(n5113) );
  INVX1 U4859 ( .A(n5074), .Y(n5121) );
  INVX1 U4860 ( .A(n5075), .Y(n5129) );
  INVX1 U4861 ( .A(n5076), .Y(n5137) );
  INVX1 U4862 ( .A(n5077), .Y(n5165) );
  INVX1 U4863 ( .A(n5078), .Y(n5173) );
  INVX1 U4864 ( .A(n5098), .Y(n5094) );
  INVX1 U4865 ( .A(n5108), .Y(n5104) );
  INVX1 U4866 ( .A(n5150), .Y(n5146) );
  INVX1 U4867 ( .A(n938), .Y(n5157) );
  INVX1 U4868 ( .A(n5073), .Y(n5114) );
  INVX1 U4869 ( .A(n5074), .Y(n5122) );
  INVX1 U4870 ( .A(n5075), .Y(n5130) );
  INVX1 U4871 ( .A(n943), .Y(n5138) );
  INVX1 U4872 ( .A(n5077), .Y(n5166) );
  INVX1 U4873 ( .A(n5078), .Y(n5174) );
  INVX1 U4874 ( .A(n5098), .Y(n5095) );
  INVX1 U4875 ( .A(n5108), .Y(n5105) );
  INVX1 U4876 ( .A(n5150), .Y(n5147) );
  INVX1 U4877 ( .A(n938), .Y(n5158) );
  INVX1 U4878 ( .A(n5073), .Y(n5115) );
  INVX1 U4879 ( .A(n5074), .Y(n5123) );
  INVX1 U4880 ( .A(n5075), .Y(n5131) );
  INVX1 U4881 ( .A(n5076), .Y(n5139) );
  INVX1 U4882 ( .A(n5077), .Y(n5167) );
  INVX1 U4883 ( .A(n5078), .Y(n5175) );
  INVX1 U4884 ( .A(n5098), .Y(n5096) );
  INVX1 U4885 ( .A(n5108), .Y(n5106) );
  INVX1 U4886 ( .A(n5150), .Y(n5148) );
  INVX1 U4887 ( .A(n5160), .Y(n5159) );
  INVX1 U4888 ( .A(n957), .Y(n5093) );
  INVX1 U4889 ( .A(n952), .Y(n5103) );
  INVX1 U4890 ( .A(n5073), .Y(n5112) );
  INVX1 U4891 ( .A(n5074), .Y(n5120) );
  INVX1 U4892 ( .A(n5075), .Y(n5128) );
  INVX1 U4893 ( .A(n5076), .Y(n5136) );
  INVX1 U4894 ( .A(n941), .Y(n5145) );
  INVX1 U4895 ( .A(n5160), .Y(n5156) );
  INVX1 U4896 ( .A(n5077), .Y(n5164) );
  INVX1 U4897 ( .A(n5078), .Y(n5172) );
  INVX1 U4898 ( .A(n5379), .Y(n5364) );
  INVX1 U4899 ( .A(n5401), .Y(n5386) );
  INVX1 U4900 ( .A(n5379), .Y(n5365) );
  INVX1 U4901 ( .A(n5401), .Y(n5387) );
  INVX1 U4902 ( .A(n5379), .Y(n5363) );
  INVX1 U4903 ( .A(n5401), .Y(n5385) );
  INVX1 U4904 ( .A(n5073), .Y(n5116) );
  INVX1 U4905 ( .A(n5074), .Y(n5124) );
  INVX1 U4906 ( .A(n5075), .Y(n5132) );
  INVX1 U4907 ( .A(n5076), .Y(n5140) );
  INVX1 U4908 ( .A(n5077), .Y(n5168) );
  INVX1 U4909 ( .A(n5078), .Y(n5176) );
  INVX1 U4910 ( .A(n5372), .Y(n5367) );
  INVX1 U4911 ( .A(n5394), .Y(n5389) );
  INVX1 U4912 ( .A(n5098), .Y(n5097) );
  INVX1 U4913 ( .A(n5108), .Y(n5107) );
  INVX1 U4914 ( .A(n5150), .Y(n5149) );
  CLKINVX3 U4915 ( .A(n5587), .Y(n5582) );
  CLKINVX3 U4916 ( .A(n5586), .Y(n5585) );
  CLKINVX3 U4917 ( .A(n5586), .Y(n5583) );
  CLKINVX3 U4918 ( .A(n5586), .Y(n5584) );
  INVX1 U4919 ( .A(n926), .Y(n5179) );
  INVX1 U4920 ( .A(n5182), .Y(n5178) );
  INVX1 U4921 ( .A(n5182), .Y(n5177) );
  INVX1 U4922 ( .A(n5182), .Y(n5181) );
  INVX1 U4923 ( .A(n5182), .Y(n5180) );
  CLKINVX3 U4924 ( .A(n5274), .Y(n5261) );
  CLKINVX3 U4925 ( .A(n5273), .Y(n5262) );
  CLKINVX3 U4926 ( .A(n5274), .Y(n5263) );
  CLKINVX3 U4927 ( .A(n5273), .Y(n5264) );
  CLKINVX3 U4928 ( .A(n5557), .Y(n5553) );
  CLKINVX3 U4929 ( .A(n5556), .Y(n5554) );
  CLKINVX3 U4930 ( .A(n5556), .Y(n5555) );
  CLKINVX3 U4931 ( .A(n5557), .Y(n5552) );
  INVX1 U4932 ( .A(n5216), .Y(n5215) );
  INVX1 U4933 ( .A(n5248), .Y(n5247) );
  INVX1 U4934 ( .A(n5216), .Y(n5214) );
  INVX1 U4935 ( .A(n5248), .Y(n5246) );
  INVX1 U4936 ( .A(n5216), .Y(n5213) );
  INVX1 U4937 ( .A(n5248), .Y(n5245) );
  CLKINVX3 U4938 ( .A(n5337), .Y(n5336) );
  CLKINVX3 U4939 ( .A(n5350), .Y(n5349) );
  CLKINVX3 U4940 ( .A(n5337), .Y(n5335) );
  CLKINVX3 U4941 ( .A(n5350), .Y(n5348) );
  CLKINVX3 U4942 ( .A(n5338), .Y(n5334) );
  CLKINVX3 U4943 ( .A(n5351), .Y(n5347) );
  INVX1 U4944 ( .A(n5074), .Y(n5117) );
  INVX1 U4945 ( .A(n5078), .Y(n5169) );
  INVX1 U4946 ( .A(n5073), .Y(n5109) );
  INVX1 U4947 ( .A(n5075), .Y(n5125) );
  INVX1 U4948 ( .A(n920), .Y(n5424) );
  INVX1 U4949 ( .A(n918), .Y(n5446) );
  INVX1 U4950 ( .A(n920), .Y(n5425) );
  INVX1 U4951 ( .A(n918), .Y(n5447) );
  INVX1 U4952 ( .A(n920), .Y(n5423) );
  INVX1 U4953 ( .A(n918), .Y(n5445) );
  INVX1 U4954 ( .A(n5801), .Y(n5150) );
  INVX1 U4955 ( .A(n913), .Y(n5500) );
  INVX1 U4956 ( .A(n911), .Y(n5522) );
  INVX1 U4957 ( .A(n913), .Y(n5501) );
  INVX1 U4958 ( .A(n911), .Y(n5523) );
  INVX1 U4959 ( .A(n913), .Y(n5502) );
  INVX1 U4960 ( .A(n911), .Y(n5524) );
  INVX1 U4961 ( .A(n5799), .Y(n5098) );
  INVX1 U4962 ( .A(n5800), .Y(n5108) );
  INVX1 U4963 ( .A(n5160), .Y(n5151) );
  INVX1 U4964 ( .A(n5802), .Y(n5160) );
  INVX1 U4965 ( .A(n917), .Y(n5456) );
  INVX1 U4966 ( .A(n915), .Y(n5478) );
  INVX1 U4967 ( .A(n917), .Y(n5457) );
  INVX1 U4968 ( .A(n915), .Y(n5479) );
  INVX1 U4969 ( .A(n916), .Y(n5467) );
  INVX1 U4970 ( .A(n914), .Y(n5489) );
  INVX1 U4971 ( .A(n909), .Y(n5544) );
  INVX1 U4972 ( .A(n887), .Y(n5579) );
  INVX1 U4973 ( .A(n916), .Y(n5468) );
  INVX1 U4974 ( .A(n914), .Y(n5490) );
  INVX1 U4975 ( .A(n909), .Y(n5545) );
  INVX1 U4976 ( .A(n887), .Y(n5580) );
  INVX1 U4977 ( .A(n921), .Y(n5414) );
  INVX1 U4978 ( .A(n919), .Y(n5436) );
  INVX1 U4979 ( .A(n921), .Y(n5413) );
  INVX1 U4980 ( .A(n919), .Y(n5435) );
  INVX1 U4981 ( .A(n921), .Y(n5412) );
  INVX1 U4982 ( .A(n919), .Y(n5434) );
  INVX1 U4983 ( .A(n912), .Y(n5513) );
  INVX1 U4984 ( .A(n910), .Y(n5535) );
  INVX1 U4985 ( .A(n912), .Y(n5512) );
  INVX1 U4986 ( .A(n910), .Y(n5534) );
  INVX1 U4987 ( .A(n912), .Y(n5511) );
  INVX1 U4988 ( .A(n910), .Y(n5533) );
  INVX1 U4989 ( .A(n5077), .Y(n5161) );
  INVX1 U4990 ( .A(n916), .Y(n5469) );
  INVX1 U4991 ( .A(n914), .Y(n5491) );
  INVX1 U4992 ( .A(n909), .Y(n5546) );
  INVX1 U4993 ( .A(n887), .Y(n5581) );
  CLKINVX3 U4994 ( .A(n5458), .Y(n5448) );
  INVX1 U4995 ( .A(n917), .Y(n5458) );
  CLKINVX3 U4996 ( .A(n5480), .Y(n5470) );
  INVX1 U4997 ( .A(n915), .Y(n5480) );
  CLKINVX3 U4998 ( .A(n5568), .Y(n5564) );
  CLKINVX3 U4999 ( .A(n5567), .Y(n5565) );
  CLKINVX3 U5000 ( .A(n5567), .Y(n5566) );
  INVX1 U5001 ( .A(n5380), .Y(n5378) );
  INVX1 U5002 ( .A(n5402), .Y(n5400) );
  CLKINVX3 U5003 ( .A(n5563), .Y(n5561) );
  INVX1 U5004 ( .A(n5563), .Y(n5562) );
  CLKINVX3 U5005 ( .A(n5593), .Y(n5588) );
  CLKINVX3 U5006 ( .A(n5592), .Y(n5589) );
  CLKINVX3 U5007 ( .A(n5592), .Y(n5590) );
  CLKINVX3 U5008 ( .A(n5592), .Y(n5591) );
  INVX1 U5009 ( .A(n922), .Y(n5185) );
  INVX1 U5010 ( .A(n5551), .Y(n5548) );
  INVX1 U5011 ( .A(n5188), .Y(n5183) );
  INVX1 U5012 ( .A(n5188), .Y(n5184) );
  INVX1 U5013 ( .A(n5551), .Y(n5547) );
  INVX1 U5014 ( .A(n5188), .Y(n5186) );
  INVX1 U5015 ( .A(n5188), .Y(n5187) );
  INVX1 U5016 ( .A(n5551), .Y(n5550) );
  INVX1 U5017 ( .A(n5551), .Y(n5549) );
  INVX1 U5018 ( .A(n5179), .Y(n5182) );
  INVX1 U5019 ( .A(n886), .Y(n5587) );
  INVX1 U5020 ( .A(n886), .Y(n5586) );
  INVX1 U5021 ( .A(n5381), .Y(n5377) );
  INVX1 U5022 ( .A(n5403), .Y(n5399) );
  INVX1 U5023 ( .A(n5380), .Y(n5376) );
  INVX1 U5024 ( .A(n5402), .Y(n5398) );
  INVX1 U5025 ( .A(n5381), .Y(n5375) );
  INVX1 U5026 ( .A(n5403), .Y(n5397) );
  INVX1 U5027 ( .A(n5381), .Y(n5374) );
  INVX1 U5028 ( .A(n5403), .Y(n5396) );
  INVX1 U5029 ( .A(n5381), .Y(n5373) );
  INVX1 U5030 ( .A(n5403), .Y(n5395) );
  INVX1 U5031 ( .A(n5381), .Y(n5372) );
  INVX1 U5032 ( .A(n5403), .Y(n5394) );
  INVX1 U5033 ( .A(n5381), .Y(n5371) );
  INVX1 U5034 ( .A(n5403), .Y(n5393) );
  INVX1 U5035 ( .A(n5380), .Y(n5370) );
  INVX1 U5036 ( .A(n5402), .Y(n5392) );
  INVX1 U5037 ( .A(n5380), .Y(n5369) );
  INVX1 U5038 ( .A(n5402), .Y(n5391) );
  INVX1 U5039 ( .A(n5381), .Y(n5368) );
  INVX1 U5040 ( .A(n5403), .Y(n5390) );
  CLKINVX3 U5041 ( .A(n5563), .Y(n5560) );
  INVX1 U5042 ( .A(n907), .Y(n5556) );
  CLKINVX3 U5043 ( .A(n5288), .Y(n5284) );
  CLKINVX3 U5044 ( .A(n5288), .Y(n5287) );
  CLKINVX3 U5045 ( .A(n5289), .Y(n5285) );
  CLKINVX3 U5046 ( .A(n5260), .Y(n5259) );
  INVX1 U5047 ( .A(n5278), .Y(n5273) );
  INVX1 U5048 ( .A(n5278), .Y(n5274) );
  INVX1 U5049 ( .A(n5280), .Y(n5265) );
  INVX1 U5050 ( .A(n5279), .Y(n5270) );
  INVX1 U5051 ( .A(n5280), .Y(n5266) );
  INVX1 U5052 ( .A(n5280), .Y(n5271) );
  INVX1 U5053 ( .A(n5279), .Y(n5269) );
  INVX1 U5054 ( .A(n5278), .Y(n5272) );
  INVX1 U5055 ( .A(n5280), .Y(n5268) );
  INVX1 U5056 ( .A(n5279), .Y(n5267) );
  CLKINVX3 U5057 ( .A(n4475), .Y(n5594) );
  CLKINVX3 U5058 ( .A(n4476), .Y(n5597) );
  CLKINVX3 U5059 ( .A(n4477), .Y(n5600) );
  CLKINVX3 U5060 ( .A(n4478), .Y(n5603) );
  CLKINVX3 U5061 ( .A(n4479), .Y(n5606) );
  CLKINVX3 U5062 ( .A(n4480), .Y(n5609) );
  CLKINVX3 U5063 ( .A(n4481), .Y(n5612) );
  CLKINVX3 U5064 ( .A(n4482), .Y(n5615) );
  CLKINVX3 U5065 ( .A(n4483), .Y(n5618) );
  CLKINVX3 U5066 ( .A(n4484), .Y(n5621) );
  CLKINVX3 U5067 ( .A(n4485), .Y(n5624) );
  CLKINVX3 U5068 ( .A(n4486), .Y(n5627) );
  CLKINVX3 U5069 ( .A(n4487), .Y(n5630) );
  CLKINVX3 U5070 ( .A(n4488), .Y(n5633) );
  CLKINVX3 U5071 ( .A(n4475), .Y(n5595) );
  CLKINVX3 U5072 ( .A(n4476), .Y(n5598) );
  CLKINVX3 U5073 ( .A(n4478), .Y(n5604) );
  CLKINVX3 U5074 ( .A(n4479), .Y(n5607) );
  CLKINVX3 U5075 ( .A(n4480), .Y(n5610) );
  CLKINVX3 U5076 ( .A(n4481), .Y(n5613) );
  CLKINVX3 U5077 ( .A(n4482), .Y(n5616) );
  CLKINVX3 U5078 ( .A(n4483), .Y(n5619) );
  CLKINVX3 U5079 ( .A(n4484), .Y(n5622) );
  CLKINVX3 U5080 ( .A(n4485), .Y(n5625) );
  CLKINVX3 U5081 ( .A(n4486), .Y(n5628) );
  CLKINVX3 U5082 ( .A(n4487), .Y(n5631) );
  CLKINVX3 U5083 ( .A(n4475), .Y(n5596) );
  CLKINVX3 U5084 ( .A(n4476), .Y(n5599) );
  CLKINVX3 U5085 ( .A(n4477), .Y(n5602) );
  CLKINVX3 U5086 ( .A(n4478), .Y(n5605) );
  CLKINVX3 U5087 ( .A(n4479), .Y(n5608) );
  CLKINVX3 U5088 ( .A(n4480), .Y(n5611) );
  CLKINVX3 U5089 ( .A(n4481), .Y(n5614) );
  CLKINVX3 U5090 ( .A(n4482), .Y(n5617) );
  CLKINVX3 U5091 ( .A(n4483), .Y(n5620) );
  CLKINVX3 U5092 ( .A(n4484), .Y(n5623) );
  CLKINVX3 U5093 ( .A(n4485), .Y(n5626) );
  CLKINVX3 U5094 ( .A(n4486), .Y(n5629) );
  CLKINVX3 U5095 ( .A(n4487), .Y(n5632) );
  CLKINVX3 U5096 ( .A(n4488), .Y(n5634) );
  CLKINVX3 U5097 ( .A(n4477), .Y(n5601) );
  CLKINVX3 U5098 ( .A(n5638), .Y(n5637) );
  CLKINVX3 U5099 ( .A(n5638), .Y(n5636) );
  CLKINVX3 U5100 ( .A(n5260), .Y(n5258) );
  CLKINVX3 U5101 ( .A(n5252), .Y(n5251) );
  INVX1 U5102 ( .A(n4488), .Y(n5635) );
  INVX1 U5103 ( .A(n5192), .Y(n5191) );
  INVX1 U5104 ( .A(n5196), .Y(n5195) );
  INVX1 U5105 ( .A(n5200), .Y(n5199) );
  INVX1 U5106 ( .A(n5204), .Y(n5203) );
  INVX1 U5107 ( .A(n5208), .Y(n5207) );
  INVX1 U5108 ( .A(n5212), .Y(n5211) );
  INVX1 U5109 ( .A(n5220), .Y(n5219) );
  INVX1 U5110 ( .A(n5224), .Y(n5223) );
  INVX1 U5111 ( .A(n5228), .Y(n5227) );
  INVX1 U5112 ( .A(n5232), .Y(n5231) );
  INVX1 U5113 ( .A(n5236), .Y(n5235) );
  INVX1 U5114 ( .A(n5240), .Y(n5239) );
  INVX1 U5115 ( .A(n5244), .Y(n5242) );
  INVX1 U5116 ( .A(n5192), .Y(n5190) );
  INVX1 U5117 ( .A(n5196), .Y(n5194) );
  INVX1 U5118 ( .A(n5200), .Y(n5198) );
  INVX1 U5119 ( .A(n5204), .Y(n5202) );
  INVX1 U5120 ( .A(n5208), .Y(n5206) );
  INVX1 U5121 ( .A(n5212), .Y(n5210) );
  INVX1 U5122 ( .A(n5220), .Y(n5218) );
  INVX1 U5123 ( .A(n5224), .Y(n5222) );
  INVX1 U5124 ( .A(n5228), .Y(n5226) );
  INVX1 U5125 ( .A(n5232), .Y(n5230) );
  INVX1 U5126 ( .A(n5236), .Y(n5234) );
  INVX1 U5127 ( .A(n5240), .Y(n5238) );
  INVX1 U5128 ( .A(n5244), .Y(n5241) );
  INVX1 U5129 ( .A(n5192), .Y(n5189) );
  INVX1 U5130 ( .A(n5196), .Y(n5193) );
  INVX1 U5131 ( .A(n5204), .Y(n5201) );
  INVX1 U5132 ( .A(n5208), .Y(n5205) );
  INVX1 U5133 ( .A(n5212), .Y(n5209) );
  INVX1 U5134 ( .A(n5220), .Y(n5217) );
  INVX1 U5135 ( .A(n5224), .Y(n5221) );
  INVX1 U5136 ( .A(n5228), .Y(n5225) );
  INVX1 U5137 ( .A(n5232), .Y(n5229) );
  INVX1 U5138 ( .A(n5236), .Y(n5233) );
  INVX1 U5139 ( .A(n5240), .Y(n5237) );
  INVX1 U5140 ( .A(n5200), .Y(n5197) );
  INVX1 U5141 ( .A(n5849), .Y(n5216) );
  INVX1 U5142 ( .A(n5857), .Y(n5248) );
  INVX1 U5143 ( .A(n5244), .Y(n5243) );
  INVX1 U5144 ( .A(n907), .Y(n5557) );
  INVX1 U5145 ( .A(n889), .Y(n5567) );
  INVX1 U5146 ( .A(n889), .Y(n5568) );
  INVX1 U5147 ( .A(n5071), .Y(n5338) );
  INVX1 U5148 ( .A(n5072), .Y(n5351) );
  INVX1 U5149 ( .A(n906), .Y(n5563) );
  NAND2X1 U5150 ( .A(n5249), .B(n926), .Y(n886) );
  INVX1 U5151 ( .A(n5185), .Y(n5188) );
  INVX1 U5152 ( .A(n885), .Y(n5593) );
  INVX1 U5153 ( .A(n885), .Y(n5592) );
  INVX1 U5154 ( .A(n908), .Y(n5551) );
  INVX1 U5155 ( .A(n942), .Y(n5380) );
  INVX1 U5156 ( .A(n940), .Y(n5402) );
  INVX1 U5157 ( .A(n942), .Y(n5381) );
  INVX1 U5158 ( .A(n940), .Y(n5403) );
  INVX1 U5159 ( .A(n5071), .Y(n5341) );
  INVX1 U5160 ( .A(n5072), .Y(n5354) );
  INVX1 U5161 ( .A(n5071), .Y(n5342) );
  INVX1 U5162 ( .A(n5072), .Y(n5355) );
  INVX1 U5163 ( .A(n5071), .Y(n5343) );
  INVX1 U5164 ( .A(n5072), .Y(n5356) );
  INVX1 U5165 ( .A(n5071), .Y(n5344) );
  INVX1 U5166 ( .A(n5072), .Y(n5357) );
  INVX1 U5167 ( .A(n5071), .Y(n5345) );
  INVX1 U5168 ( .A(n5072), .Y(n5358) );
  INVX1 U5169 ( .A(n5071), .Y(n5346) );
  INVX1 U5170 ( .A(n5072), .Y(n5359) );
  INVX1 U5171 ( .A(n5071), .Y(n5339) );
  INVX1 U5172 ( .A(n5072), .Y(n5352) );
  INVX1 U5173 ( .A(n5071), .Y(n5340) );
  INVX1 U5174 ( .A(n5072), .Y(n5353) );
  NAND2X1 U5175 ( .A(n932), .B(n5250), .Y(n907) );
  CLKINVX3 U5176 ( .A(n4915), .Y(n4916) );
  CLKINVX3 U5177 ( .A(n4915), .Y(n4917) );
  CLKINVX3 U5178 ( .A(n4905), .Y(n4906) );
  CLKINVX3 U5179 ( .A(n4920), .Y(n4921) );
  CLKINVX3 U5180 ( .A(n4909), .Y(n4910) );
  CLKINVX3 U5181 ( .A(n4897), .Y(n4898) );
  CLKINVX3 U5182 ( .A(n4901), .Y(n4902) );
  CLKINVX3 U5183 ( .A(n4893), .Y(n4894) );
  CLKINVX3 U5184 ( .A(n4913), .Y(n4914) );
  CLKINVX3 U5185 ( .A(n4903), .Y(n4904) );
  CLKINVX3 U5186 ( .A(n4918), .Y(n4919) );
  CLKINVX3 U5187 ( .A(n4907), .Y(n4908) );
  CLKINVX3 U5188 ( .A(n4895), .Y(n4896) );
  CLKINVX3 U5189 ( .A(n4899), .Y(n4900) );
  CLKINVX3 U5190 ( .A(n4891), .Y(n4892) );
  CLKINVX3 U5191 ( .A(n4911), .Y(n4912) );
  CLKINVX3 U5192 ( .A(n5313), .Y(n5305) );
  CLKINVX3 U5193 ( .A(n5312), .Y(n5306) );
  CLKINVX3 U5194 ( .A(n5312), .Y(n5307) );
  CLKINVX3 U5195 ( .A(n5295), .Y(n5286) );
  CLKINVX3 U5196 ( .A(n5311), .Y(n5309) );
  CLKINVX3 U5197 ( .A(n5311), .Y(n5308) );
  CLKINVX3 U5198 ( .A(n5311), .Y(n5310) );
  INVX4 U5199 ( .A(n5300), .Y(n5299) );
  CLKINVX3 U5200 ( .A(n5322), .Y(n5317) );
  CLKINVX3 U5201 ( .A(n5323), .Y(n5319) );
  CLKINVX3 U5202 ( .A(n5322), .Y(n5320) );
  CLKINVX3 U5203 ( .A(n5322), .Y(n5318) );
  CLKINVX3 U5204 ( .A(n5323), .Y(n5321) );
  INVX1 U5205 ( .A(n5297), .Y(n5288) );
  INVX1 U5206 ( .A(n5279), .Y(n5275) );
  INVX1 U5207 ( .A(n5280), .Y(n5276) );
  INVX1 U5208 ( .A(n5281), .Y(n5278) );
  INVX1 U5209 ( .A(n5281), .Y(n5280) );
  INVX1 U5210 ( .A(n5281), .Y(n5279) );
  INVX1 U5211 ( .A(n5279), .Y(n5277) );
  CLKINVX3 U5212 ( .A(n5328), .Y(n5327) );
  CLKINVX3 U5213 ( .A(n5256), .Y(n5253) );
  CLKINVX3 U5214 ( .A(n5301), .Y(n5298) );
  CLKINVX3 U5215 ( .A(n5303), .Y(n5302) );
  CLKINVX3 U5216 ( .A(n5260), .Y(n5257) );
  INVX1 U5217 ( .A(n1322), .Y(n5260) );
  INVX1 U5218 ( .A(n874), .Y(n5849) );
  INVX1 U5219 ( .A(n858), .Y(n5857) );
  CLKINVX3 U5220 ( .A(n5326), .Y(n5325) );
  CLKINVX3 U5221 ( .A(n5326), .Y(n5324) );
  CLKINVX3 U5222 ( .A(n5255), .Y(n5254) );
  INVX12 U5223 ( .A(n5283), .Y(n5282) );
  INVX1 U5224 ( .A(n5845), .Y(n5200) );
  INVX1 U5225 ( .A(n5853), .Y(n5232) );
  INVX1 U5226 ( .A(n5854), .Y(n5236) );
  INVX1 U5227 ( .A(n5846), .Y(n5204) );
  INVX1 U5228 ( .A(n5850), .Y(n5220) );
  INVX1 U5229 ( .A(n5855), .Y(n5240) );
  INVX1 U5230 ( .A(n5843), .Y(n5192) );
  INVX1 U5231 ( .A(n5847), .Y(n5208) );
  INVX1 U5232 ( .A(n5851), .Y(n5224) );
  INVX1 U5233 ( .A(n5856), .Y(n5244) );
  INVX1 U5234 ( .A(n5844), .Y(n5196) );
  INVX1 U5235 ( .A(n5848), .Y(n5212) );
  INVX1 U5236 ( .A(n5852), .Y(n5228) );
  INVX1 U5237 ( .A(n757), .Y(n5638) );
  INVX1 U5238 ( .A(n1455), .Y(n5252) );
  INVX1 U5239 ( .A(n5297), .Y(n5291) );
  INVX1 U5240 ( .A(n5286), .Y(n5292) );
  INVX1 U5241 ( .A(n5297), .Y(n5293) );
  INVX1 U5242 ( .A(n5297), .Y(n5294) );
  INVX1 U5243 ( .A(n5297), .Y(n5289) );
  INVX1 U5244 ( .A(n5286), .Y(n5290) );
  INVX1 U5245 ( .A(n5297), .Y(n5295) );
  INVX1 U5246 ( .A(n5297), .Y(n5296) );
  NAND2X1 U5247 ( .A(n931), .B(n906), .Y(n889) );
  BUFX3 U5248 ( .A(n947), .Y(n5073) );
  OAI31X1 U5249 ( .A0(n944), .A1(n5859), .A2(n935), .B0(n925), .Y(n947) );
  BUFX3 U5250 ( .A(n945), .Y(n5075) );
  OAI31X1 U5251 ( .A0(n944), .A1(n5859), .A2(n930), .B0(n925), .Y(n945) );
  BUFX3 U5252 ( .A(n946), .Y(n5074) );
  OAI31X1 U5253 ( .A0(n944), .A1(n5859), .A2(n933), .B0(n925), .Y(n946) );
  BUFX3 U5254 ( .A(n943), .Y(n5076) );
  OAI31X1 U5255 ( .A0(n944), .A1(n927), .A2(n5859), .B0(n925), .Y(n943) );
  BUFX3 U5256 ( .A(n934), .Y(n5077) );
  OAI31X1 U5257 ( .A0(n935), .A1(n928), .A2(n5859), .B0(n925), .Y(n934) );
  BUFX3 U5258 ( .A(n929), .Y(n5078) );
  OAI31X1 U5259 ( .A0(n930), .A1(n928), .A2(n5859), .B0(n925), .Y(n929) );
  BUFX3 U5260 ( .A(n954), .Y(n5071) );
  OAI31X1 U5261 ( .A0(n949), .A1(n5859), .A2(n933), .B0(n925), .Y(n954) );
  BUFX3 U5262 ( .A(n948), .Y(n5072) );
  OAI31X1 U5263 ( .A0(n949), .A1(n927), .A2(n5859), .B0(n925), .Y(n948) );
  INVX1 U5264 ( .A(n925), .Y(n5797) );
  NAND2X1 U5265 ( .A(n5249), .B(n922), .Y(n885) );
  BUFX3 U5266 ( .A(n1096), .Y(n5069) );
  NOR3X1 U5267 ( .A(n5822), .B(n5823), .C(n5821), .Y(n1096) );
  INVX4 U5268 ( .A(n5332), .Y(n5330) );
  CLKINVX3 U5269 ( .A(n5332), .Y(n5331) );
  CLKINVX3 U5270 ( .A(n1128), .Y(n5885) );
  NAND2X1 U5271 ( .A(n950), .B(n5880), .Y(n933) );
  INVX8 U5272 ( .A(n4491), .Y(n5569) );
  INVX1 U5273 ( .A(n5065), .Y(n5860) );
  INVX1 U5274 ( .A(n4882), .Y(n4915) );
  INVX1 U5275 ( .A(n4884), .Y(n4920) );
  INVX1 U5276 ( .A(n4871), .Y(n4901) );
  INVX1 U5277 ( .A(n4867), .Y(n4893) );
  INVX1 U5278 ( .A(n4873), .Y(n4905) );
  INVX1 U5279 ( .A(n4869), .Y(n4897) );
  INVX1 U5280 ( .A(n4879), .Y(n4909) );
  INVX1 U5281 ( .A(n4872), .Y(n4903) );
  INVX1 U5282 ( .A(n4868), .Y(n4895) );
  INVX1 U5283 ( .A(n4878), .Y(n4907) );
  INVX1 U5284 ( .A(n4880), .Y(n4911) );
  INVX1 U5285 ( .A(n4881), .Y(n4913) );
  INVX1 U5286 ( .A(n4883), .Y(n4918) );
  INVX1 U5287 ( .A(n4870), .Y(n4899) );
  INVX1 U5288 ( .A(n4866), .Y(n4891) );
  CLKINVX3 U5289 ( .A(n931), .Y(n5859) );
  AND2X2 U5290 ( .A(n1318), .B(n5894), .Y(n1322) );
  OR2X2 U5291 ( .A(n927), .B(n928), .Y(n924) );
  CLKINVX3 U5292 ( .A(n5313), .Y(n5304) );
  INVX1 U5293 ( .A(n1185), .Y(n5313) );
  NAND2X1 U5294 ( .A(n5881), .B(n5882), .Y(n949) );
  NAND2X1 U5295 ( .A(n953), .B(n5880), .Y(n935) );
  INVX1 U5296 ( .A(n1185), .Y(n5311) );
  INVX1 U5297 ( .A(n1185), .Y(n5312) );
  INVX1 U5298 ( .A(n1189), .Y(n5300) );
  INVX1 U5299 ( .A(n1182), .Y(n5322) );
  CLKINVX3 U5300 ( .A(n5323), .Y(n5316) );
  INVX1 U5301 ( .A(n1182), .Y(n5323) );
  INVX1 U5302 ( .A(n1257), .Y(n5281) );
  BUFX3 U5303 ( .A(n1186), .Y(n5060) );
  NOR2X1 U5304 ( .A(n5894), .B(n5057), .Y(n1186) );
  INVX1 U5305 ( .A(n755), .Y(n5972) );
  NAND2X1 U5306 ( .A(n5050), .B(n858), .Y(n757) );
  BUFX3 U5307 ( .A(n1588), .Y(n5059) );
  AND2X2 U5308 ( .A(n5053), .B(n5894), .Y(n1588) );
  INVX1 U5309 ( .A(n883), .Y(n5844) );
  INVX1 U5310 ( .A(n876), .Y(n5848) );
  INVX1 U5311 ( .A(n870), .Y(n5852) );
  INVX1 U5312 ( .A(n861), .Y(n5856) );
  INVX1 U5313 ( .A(n884), .Y(n5843) );
  INVX1 U5314 ( .A(n877), .Y(n5847) );
  INVX1 U5315 ( .A(n871), .Y(n5851) );
  INVX1 U5316 ( .A(n878), .Y(n5846) );
  INVX1 U5317 ( .A(n872), .Y(n5850) );
  INVX1 U5318 ( .A(n863), .Y(n5855) );
  INVX1 U5319 ( .A(n868), .Y(n5853) );
  INVX1 U5320 ( .A(n865), .Y(n5854) );
  INVX1 U5321 ( .A(n880), .Y(n5845) );
  BUFX3 U5322 ( .A(n5877), .Y(n5051) );
  BUFX3 U5323 ( .A(n5877), .Y(n5052) );
  AND2X2 U5324 ( .A(n5055), .B(n5894), .Y(n1455) );
  INVX1 U5325 ( .A(n1139), .Y(n5326) );
  INVX1 U5326 ( .A(n1389), .Y(n5255) );
  INVX1 U5327 ( .A(n1389), .Y(n5256) );
  INVX1 U5328 ( .A(n1189), .Y(n5301) );
  INVX1 U5329 ( .A(n1188), .Y(n5303) );
  INVX1 U5330 ( .A(n1183), .Y(n5315) );
  INVX1 U5331 ( .A(n1138), .Y(n5328) );
  INVX1 U5332 ( .A(n1255), .Y(n5283) );
  CLKINVX3 U5333 ( .A(n4491), .Y(n5570) );
  INVX1 U5334 ( .A(n1254), .Y(n5297) );
  CLKINVX3 U5335 ( .A(ns[2]), .Y(n5823) );
  NOR2X2 U5336 ( .A(n960), .B(n5797), .Y(n961) );
  OAI21XL U5337 ( .A0(n923), .A1(n924), .B0(n925), .Y(n922) );
  OR3XL U5338 ( .A(ns[0]), .B(ns[1]), .C(n5823), .Y(n4490) );
  INVX1 U5339 ( .A(n1111), .Y(n5805) );
  AOI22X1 U5340 ( .A0(N1304), .A1(n4474), .B0(in_start_addr[2]), .B1(n5069), 
        .Y(n1111) );
  INVX1 U5341 ( .A(n1102), .Y(n5814) );
  AOI22X1 U5342 ( .A0(N1332), .A1(n4474), .B0(weight_start_addr[2]), .B1(n5069), .Y(n1102) );
  INVX1 U5343 ( .A(n1106), .Y(n5810) );
  AOI22X1 U5344 ( .A0(N1309), .A1(n4473), .B0(in_start_addr[7]), .B1(n5069), 
        .Y(n1106) );
  INVX1 U5345 ( .A(n1107), .Y(n5809) );
  AOI22X1 U5346 ( .A0(N1308), .A1(n4473), .B0(in_start_addr[6]), .B1(n5069), 
        .Y(n1107) );
  INVX1 U5347 ( .A(n1097), .Y(n5819) );
  AOI22X1 U5348 ( .A0(N1337), .A1(n5068), .B0(weight_start_addr[7]), .B1(n5069), .Y(n1097) );
  INVX1 U5349 ( .A(n4490), .Y(n5068) );
  INVX1 U5350 ( .A(n1098), .Y(n5818) );
  AOI22X1 U5351 ( .A0(N1336), .A1(n5067), .B0(weight_start_addr[6]), .B1(n5069), .Y(n1098) );
  INVX1 U5352 ( .A(n4490), .Y(n5067) );
  INVX1 U5353 ( .A(n1112), .Y(n5804) );
  AOI22X1 U5354 ( .A0(N1303), .A1(n5068), .B0(in_start_addr[1]), .B1(n5069), 
        .Y(n1112) );
  INVX1 U5355 ( .A(n1105), .Y(n5811) );
  AOI22X1 U5356 ( .A0(N1310), .A1(n4473), .B0(in_start_addr[8]), .B1(n5069), 
        .Y(n1105) );
  INVX1 U5357 ( .A(n1108), .Y(n5808) );
  AOI22X1 U5358 ( .A0(N1307), .A1(n4473), .B0(in_start_addr[5]), .B1(n5069), 
        .Y(n1108) );
  INVX1 U5359 ( .A(n1109), .Y(n5807) );
  AOI22X1 U5360 ( .A0(N1306), .A1(n4473), .B0(in_start_addr[4]), .B1(n5069), 
        .Y(n1109) );
  INVX1 U5361 ( .A(n1110), .Y(n5806) );
  AOI22X1 U5362 ( .A0(N1305), .A1(n5068), .B0(in_start_addr[3]), .B1(n5069), 
        .Y(n1110) );
  INVX1 U5363 ( .A(n1095), .Y(n5820) );
  AOI22X1 U5364 ( .A0(N1338), .A1(n5067), .B0(weight_start_addr[8]), .B1(n5069), .Y(n1095) );
  INVX1 U5365 ( .A(n1099), .Y(n5817) );
  AOI22X1 U5366 ( .A0(N1335), .A1(n5068), .B0(weight_start_addr[5]), .B1(n5069), .Y(n1099) );
  INVX1 U5367 ( .A(n1100), .Y(n5816) );
  AOI22X1 U5368 ( .A0(N1334), .A1(n4474), .B0(weight_start_addr[4]), .B1(n5069), .Y(n1100) );
  INVX1 U5369 ( .A(n1101), .Y(n5815) );
  AOI22X1 U5370 ( .A0(N1333), .A1(n4473), .B0(weight_start_addr[3]), .B1(n5069), .Y(n1101) );
  INVX1 U5371 ( .A(n1103), .Y(n5813) );
  AOI22X1 U5372 ( .A0(N1331), .A1(n4474), .B0(weight_start_addr[1]), .B1(n5069), .Y(n1103) );
  NOR3X1 U5373 ( .A(ns[1]), .B(ns[2]), .C(n5821), .Y(n1011) );
  OAI2BB1X1 U5374 ( .A0N(N12244), .A1N(n1136), .B0(n1140), .Y(N12604) );
  AOI22X1 U5375 ( .A0(N12124), .A1(n5327), .B0(N12524), .B1(n5325), .Y(n1140)
         );
  OAI2BB1X1 U5376 ( .A0N(N12243), .A1N(n5063), .B0(n1141), .Y(N12603) );
  AOI22X1 U5377 ( .A0(N12123), .A1(n5327), .B0(N12523), .B1(n5325), .Y(n1141)
         );
  OAI2BB1X1 U5378 ( .A0N(N12242), .A1N(n5062), .B0(n1142), .Y(N12602) );
  AOI22X1 U5379 ( .A0(N12122), .A1(n5327), .B0(N12522), .B1(n5325), .Y(n1142)
         );
  OAI2BB1X1 U5380 ( .A0N(N12241), .A1N(n1136), .B0(n1143), .Y(N12601) );
  AOI22X1 U5381 ( .A0(N12121), .A1(n5327), .B0(N12521), .B1(n5325), .Y(n1143)
         );
  INVX1 U5382 ( .A(n970), .Y(n5332) );
  CLKINVX3 U5383 ( .A(n5333), .Y(n5329) );
  INVX1 U5384 ( .A(n970), .Y(n5333) );
  CLKINVX3 U5385 ( .A(n1002), .Y(n5832) );
  OAI2BB1X1 U5386 ( .A0N(N12237), .A1N(n5063), .B0(n1147), .Y(N12597) );
  AOI22X1 U5387 ( .A0(N12117), .A1(n5327), .B0(N12517), .B1(n5325), .Y(n1147)
         );
  OAI2BB1X1 U5388 ( .A0N(N12240), .A1N(n5063), .B0(n1144), .Y(N12600) );
  AOI22X1 U5389 ( .A0(N12120), .A1(n5327), .B0(N12520), .B1(n5325), .Y(n1144)
         );
  OAI2BB1X1 U5390 ( .A0N(N12239), .A1N(n5062), .B0(n1145), .Y(N12599) );
  AOI22X1 U5391 ( .A0(N12119), .A1(n5327), .B0(N12519), .B1(n5325), .Y(n1145)
         );
  OAI2BB1X1 U5392 ( .A0N(N12238), .A1N(n1136), .B0(n1146), .Y(N12598) );
  AOI22X1 U5393 ( .A0(N12118), .A1(n5327), .B0(N12518), .B1(n5325), .Y(n1146)
         );
  OAI2BB1X1 U5394 ( .A0N(N12236), .A1N(n5062), .B0(n1148), .Y(N12596) );
  AOI22X1 U5395 ( .A0(N12116), .A1(n5327), .B0(N12516), .B1(n5325), .Y(n1148)
         );
  OAI2BB1X1 U5396 ( .A0N(N12235), .A1N(n1136), .B0(n1149), .Y(N12595) );
  AOI22X1 U5397 ( .A0(N12115), .A1(n5327), .B0(N12515), .B1(n5325), .Y(n1149)
         );
  OAI2BB1X1 U5398 ( .A0N(N12234), .A1N(n5063), .B0(n1150), .Y(N12594) );
  AOI22X1 U5399 ( .A0(N12114), .A1(n5327), .B0(N12514), .B1(n5325), .Y(n1150)
         );
  OAI2BB1X1 U5400 ( .A0N(N12233), .A1N(n5062), .B0(n1151), .Y(N12593) );
  AOI22X1 U5401 ( .A0(N12113), .A1(n5327), .B0(N12513), .B1(n5325), .Y(n1151)
         );
  OAI2BB1X1 U5402 ( .A0N(N12232), .A1N(n1136), .B0(n1152), .Y(N12592) );
  AOI22X1 U5403 ( .A0(N12112), .A1(n5327), .B0(N12512), .B1(n5325), .Y(n1152)
         );
  OAI2BB1X1 U5404 ( .A0N(N12231), .A1N(n5063), .B0(n1153), .Y(N12591) );
  AOI22X1 U5405 ( .A0(N12111), .A1(n5327), .B0(N12511), .B1(n5324), .Y(n1153)
         );
  OAI2BB1X1 U5406 ( .A0N(N12230), .A1N(n5062), .B0(n1154), .Y(N12590) );
  AOI22X1 U5407 ( .A0(N12110), .A1(n1138), .B0(N12510), .B1(n5324), .Y(n1154)
         );
  OAI2BB1X1 U5408 ( .A0N(N12229), .A1N(n1136), .B0(n1155), .Y(N12589) );
  AOI22X1 U5409 ( .A0(N12109), .A1(n5327), .B0(N12509), .B1(n5324), .Y(n1155)
         );
  OAI2BB1X1 U5410 ( .A0N(N12228), .A1N(n5063), .B0(n1156), .Y(N12588) );
  AOI22X1 U5411 ( .A0(N12108), .A1(n1138), .B0(N12508), .B1(n5324), .Y(n1156)
         );
  OAI2BB1X1 U5412 ( .A0N(N12227), .A1N(n5062), .B0(n1157), .Y(N12587) );
  AOI22X1 U5413 ( .A0(N12107), .A1(n5327), .B0(N12507), .B1(n5324), .Y(n1157)
         );
  OAI2BB1X1 U5414 ( .A0N(N12226), .A1N(n1136), .B0(n1158), .Y(N12586) );
  AOI22X1 U5415 ( .A0(N12106), .A1(n1138), .B0(N12506), .B1(n5324), .Y(n1158)
         );
  OAI2BB1X1 U5416 ( .A0N(N12225), .A1N(n5063), .B0(n1159), .Y(N12585) );
  AOI22X1 U5417 ( .A0(N12105), .A1(n1138), .B0(N12505), .B1(n5324), .Y(n1159)
         );
  OAI2BB1X1 U5418 ( .A0N(N12224), .A1N(n5062), .B0(n1160), .Y(N12584) );
  AOI22X1 U5419 ( .A0(N12104), .A1(n1138), .B0(N12504), .B1(n5324), .Y(n1160)
         );
  OAI2BB1X1 U5420 ( .A0N(N12223), .A1N(n1136), .B0(n1161), .Y(N12583) );
  AOI22X1 U5421 ( .A0(N12103), .A1(n1138), .B0(N12503), .B1(n5324), .Y(n1161)
         );
  OAI2BB1X1 U5422 ( .A0N(N12222), .A1N(n5063), .B0(n1162), .Y(N12582) );
  AOI22X1 U5423 ( .A0(N12102), .A1(n1138), .B0(N12502), .B1(n5324), .Y(n1162)
         );
  OAI2BB1X1 U5424 ( .A0N(N12221), .A1N(n5062), .B0(n1163), .Y(N12581) );
  AOI22X1 U5425 ( .A0(N12101), .A1(n1138), .B0(N12501), .B1(n5324), .Y(n1163)
         );
  CLKINVX3 U5426 ( .A(n5064), .Y(n5887) );
  AND3X2 U5427 ( .A(n5949), .B(n5950), .C(n823), .Y(n787) );
  OAI21XL U5428 ( .A0(n882), .A1(n1045), .B0(n866), .Y(n1129) );
  AND3X2 U5429 ( .A(n5954), .B(n5955), .C(n813), .Y(n835) );
  AND3X2 U5430 ( .A(n5957), .B(n5958), .C(n830), .Y(n813) );
  AND4X2 U5431 ( .A(n828), .B(n5085), .C(n5963), .D(n5964), .Y(n837) );
  AND3X2 U5432 ( .A(n5959), .B(n5960), .C(n824), .Y(n830) );
  AND3X2 U5433 ( .A(n5940), .B(n5942), .C(n822), .Y(n829) );
  AND3X2 U5434 ( .A(n5951), .B(n5952), .C(n836), .Y(n823) );
  AND2X2 U5435 ( .A(n837), .B(n5961), .Y(n824) );
  AND2X2 U5436 ( .A(n835), .B(n5953), .Y(n836) );
  AND2X2 U5437 ( .A(n854), .B(n5965), .Y(n828) );
  AND4X2 U5438 ( .A(n829), .B(n5937), .C(n5938), .D(n5939), .Y(n832) );
  AND3X2 U5439 ( .A(n5966), .B(n5967), .C(n779), .Y(n854) );
  AND2X2 U5440 ( .A(n856), .B(n5943), .Y(n822) );
  AND3X2 U5441 ( .A(n835), .B(n5944), .C(n834), .Y(n856) );
  OAI2BB1X1 U5442 ( .A0N(N12220), .A1N(n1136), .B0(n1164), .Y(N12580) );
  AOI22X1 U5443 ( .A0(N12100), .A1(n1138), .B0(N12500), .B1(n5324), .Y(n1164)
         );
  OAI2BB1X1 U5444 ( .A0N(N12219), .A1N(n5063), .B0(n1165), .Y(N12579) );
  AOI22X1 U5445 ( .A0(N12099), .A1(n1138), .B0(N12499), .B1(n5324), .Y(n1165)
         );
  OAI2BB1X1 U5446 ( .A0N(N12218), .A1N(n5062), .B0(n1166), .Y(N12578) );
  AOI22X1 U5447 ( .A0(N12098), .A1(n1138), .B0(N12498), .B1(n5324), .Y(n1166)
         );
  OAI2BB1X1 U5448 ( .A0N(N12217), .A1N(n1136), .B0(n1167), .Y(N12577) );
  AOI22X1 U5449 ( .A0(N12097), .A1(n1138), .B0(N12497), .B1(n5324), .Y(n1167)
         );
  AOI21X1 U5450 ( .A0(n1066), .A1(n1067), .B0(n5974), .Y(n1065) );
  AOI22X1 U5451 ( .A0(value_out[28]), .A1(n1059), .B0(value_out[31]), .B1(
        n1060), .Y(n1067) );
  AOI22X1 U5452 ( .A0(value_out[30]), .A1(n1061), .B0(value_out[29]), .B1(
        n1062), .Y(n1066) );
  NOR2BX1 U5453 ( .AN(n955), .B(n956), .Y(n950) );
  NAND2X1 U5454 ( .A(n936), .B(n937), .Y(n928) );
  INVX1 U5455 ( .A(n1012), .Y(n5973) );
  OR2X2 U5456 ( .A(length_out[1]), .B(length_out[0]), .Y(n5640) );
  INVX1 U5457 ( .A(n873), .Y(n5842) );
  BUFX3 U5458 ( .A(n762), .Y(n5079) );
  NOR4X1 U5459 ( .A(n821), .B(n826), .C(n838), .D(n839), .Y(n762) );
  NAND4X1 U5460 ( .A(n801), .B(n814), .C(n784), .D(n777), .Y(n839) );
  NAND2BX1 U5461 ( .AN(n833), .B(n840), .Y(n838) );
  BUFX3 U5462 ( .A(n759), .Y(n5082) );
  NOR4X1 U5463 ( .A(n795), .B(n796), .C(n797), .D(n798), .Y(n759) );
  NAND4X1 U5464 ( .A(n799), .B(n800), .C(n801), .D(n802), .Y(n798) );
  NAND3X1 U5465 ( .A(n815), .B(n5970), .C(n816), .Y(n797) );
  AND2X2 U5466 ( .A(n1059), .B(n5974), .Y(n1044) );
  BUFX3 U5467 ( .A(n860), .Y(n5065) );
  NAND3X1 U5468 ( .A(n5890), .B(n5889), .C(n1118), .Y(n860) );
  NAND2X1 U5469 ( .A(n1120), .B(n1121), .Y(n1115) );
  AOI222X1 U5470 ( .A0(value_out[1]), .A1(n1062), .B0(value_out[3]), .B1(n1060), .C0(value_out[2]), .C1(n1061), .Y(n1080) );
  AOI222X1 U5471 ( .A0(value_out[9]), .A1(n1062), .B0(value_out[11]), .B1(
        n1060), .C0(value_out[10]), .C1(n1061), .Y(n1075) );
  AOI222X1 U5472 ( .A0(value_out[17]), .A1(n1062), .B0(value_out[19]), .B1(
        n1060), .C0(value_out[18]), .C1(n1061), .Y(n1063) );
  AOI222X1 U5473 ( .A0(value_out[33]), .A1(n1062), .B0(value_out[35]), .B1(
        n1060), .C0(value_out[34]), .C1(n1061), .Y(n1085) );
  OAI2BB1X1 U5474 ( .A0N(N12216), .A1N(n5063), .B0(n1168), .Y(N12576) );
  AOI22X1 U5475 ( .A0(N12096), .A1(n1138), .B0(N12496), .B1(n5325), .Y(n1168)
         );
  OAI2BB1X1 U5476 ( .A0N(N12215), .A1N(n5062), .B0(n1169), .Y(N12575) );
  AOI22X1 U5477 ( .A0(N12095), .A1(n1138), .B0(N12495), .B1(n5324), .Y(n1169)
         );
  OAI2BB1X1 U5478 ( .A0N(N12214), .A1N(n1136), .B0(n1170), .Y(N12574) );
  AOI22X1 U5479 ( .A0(N12094), .A1(n1138), .B0(N12494), .B1(n5325), .Y(n1170)
         );
  OAI2BB1X1 U5480 ( .A0N(N12213), .A1N(n5063), .B0(n1171), .Y(N12573) );
  AOI22X1 U5481 ( .A0(N12093), .A1(n1138), .B0(N12493), .B1(n5324), .Y(n1171)
         );
  AND2X2 U5482 ( .A(mem_num_0), .B(n5250), .Y(n4491) );
  NOR3X2 U5483 ( .A(n754), .B(n5972), .C(n753), .Y(n1032) );
  AND2X2 U5484 ( .A(n753), .B(n5841), .Y(n1031) );
  NAND3X2 U5485 ( .A(n1649), .B(n5894), .C(n1648), .Y(n1656) );
  INVX1 U5486 ( .A(n937), .Y(n5881) );
  NAND2X1 U5487 ( .A(n936), .B(n5881), .Y(n939) );
  INVX1 U5488 ( .A(n936), .Y(n5882) );
  NOR3X1 U5489 ( .A(n5088), .B(n5087), .C(n5891), .Y(n1583) );
  NAND2X1 U5490 ( .A(n937), .B(n5882), .Y(n944) );
  NOR3X1 U5491 ( .A(n5892), .B(n5087), .C(n5891), .Y(n1450) );
  BUFX3 U5492 ( .A(n1250), .Y(n5057) );
  NAND3X1 U5493 ( .A(n5088), .B(n5891), .C(n5087), .Y(n1250) );
  NAND2X1 U5494 ( .A(n950), .B(n951), .Y(n927) );
  NOR2X1 U5495 ( .A(n5057), .B(n5086), .Y(n1255) );
  NAND2X1 U5496 ( .A(n953), .B(n951), .Y(n930) );
  AND2X2 U5497 ( .A(n956), .B(n955), .Y(n953) );
  INVX1 U5498 ( .A(n754), .Y(n5841) );
  OAI2BB1X1 U5499 ( .A0N(N12212), .A1N(n5062), .B0(n1172), .Y(N12572) );
  AOI22X1 U5500 ( .A0(N12092), .A1(n1138), .B0(N12492), .B1(n5325), .Y(n1172)
         );
  OAI2BB1X1 U5501 ( .A0N(N12211), .A1N(n1136), .B0(n1173), .Y(N12571) );
  AOI22X1 U5502 ( .A0(N12091), .A1(n1138), .B0(N12491), .B1(n5324), .Y(n1173)
         );
  OAI2BB1X1 U5503 ( .A0N(N12210), .A1N(n5063), .B0(n1174), .Y(N12570) );
  AOI22X1 U5504 ( .A0(N12090), .A1(n1138), .B0(N12490), .B1(n5325), .Y(n1174)
         );
  OAI2BB1X1 U5505 ( .A0N(N12209), .A1N(n5062), .B0(n1175), .Y(N12569) );
  AOI22X1 U5506 ( .A0(N12089), .A1(n1138), .B0(N12489), .B1(n1139), .Y(n1175)
         );
  AND2X2 U5507 ( .A(n5055), .B(n5086), .Y(n1189) );
  AND3X2 U5508 ( .A(n792), .B(n793), .C(n794), .Y(n789) );
  AND2X2 U5509 ( .A(N11312), .B(n1649), .Y(N11320) );
  AND2X2 U5510 ( .A(N11311), .B(n1649), .Y(N11319) );
  AND2X2 U5511 ( .A(N11310), .B(n1649), .Y(N11318) );
  AND2X2 U5512 ( .A(N11309), .B(n1649), .Y(N11317) );
  AND2X2 U5513 ( .A(N11308), .B(n1649), .Y(N11316) );
  AND2X2 U5514 ( .A(N11307), .B(n1649), .Y(N11315) );
  INVX1 U5515 ( .A(n5061), .Y(n5663) );
  AOI21X1 U5516 ( .A0(n5972), .A1(n1012), .B0(n746), .Y(n747) );
  NOR3X1 U5517 ( .A(n746), .B(n747), .C(n4890), .Y(n741) );
  AND2X2 U5518 ( .A(n5061), .B(n5050), .Y(n5062) );
  AND2X2 U5519 ( .A(n5061), .B(n5050), .Y(n1136) );
  AND2X2 U5520 ( .A(n5061), .B(n5050), .Y(n5063) );
  NOR2X1 U5521 ( .A(n753), .B(n754), .Y(n750) );
  NOR2X1 U5522 ( .A(n873), .B(n5887), .Y(n1139) );
  AOI21X1 U5523 ( .A0(n4890), .A1(n5878), .B0(n747), .Y(n743) );
  NAND3X1 U5524 ( .A(n5938), .B(n5939), .C(n5967), .Y(n847) );
  NAND3X1 U5525 ( .A(n5957), .B(n5958), .C(n5955), .Y(n849) );
  NAND3X1 U5526 ( .A(n5085), .B(n5963), .C(n5961), .Y(n848) );
  AOI21X1 U5527 ( .A0(n862), .A1(n864), .B0(n1092), .Y(N14271) );
  AND2X2 U5528 ( .A(n1384), .B(n5894), .Y(n1389) );
  BUFX3 U5529 ( .A(n756), .Y(n5084) );
  AND4X2 U5530 ( .A(n777), .B(n778), .C(n779), .D(n780), .Y(n756) );
  AND4X2 U5531 ( .A(n5085), .B(n781), .C(n782), .D(n5966), .Y(n780) );
  AND2X2 U5532 ( .A(n1318), .B(n5086), .Y(n1187) );
  AND2X2 U5533 ( .A(n1384), .B(n5086), .Y(n1188) );
  AND4X2 U5534 ( .A(n834), .B(n5942), .C(n5940), .D(n5943), .Y(n843) );
  OAI2BB1X1 U5535 ( .A0N(N12208), .A1N(n1136), .B0(n1176), .Y(N12568) );
  AOI22X1 U5536 ( .A0(N12088), .A1(n1138), .B0(N12488), .B1(n1139), .Y(n1176)
         );
  OAI2BB1X1 U5537 ( .A0N(N12207), .A1N(n5063), .B0(n1177), .Y(N12567) );
  AOI22X1 U5538 ( .A0(N12087), .A1(n1138), .B0(N12487), .B1(n1139), .Y(n1177)
         );
  AND2X2 U5539 ( .A(n5056), .B(n5894), .Y(n1522) );
  AND2X2 U5540 ( .A(n5056), .B(n5086), .Y(n1183) );
  CLKINVX3 U5541 ( .A(n5087), .Y(n5893) );
  INVX1 U5542 ( .A(n5088), .Y(n5892) );
  AND2X2 U5543 ( .A(N1356), .B(n5250), .Y(N1364) );
  AND2X2 U5544 ( .A(N1355), .B(n5250), .Y(N1363) );
  AND2X2 U5545 ( .A(N1357), .B(n5250), .Y(N1365) );
  AND2X2 U5546 ( .A(N1358), .B(n5250), .Y(N1366) );
  AND2X2 U5547 ( .A(N1360), .B(n5250), .Y(N1368) );
  AND2X2 U5548 ( .A(N1359), .B(n5250), .Y(N1367) );
  OAI2BB1X1 U5549 ( .A0N(n5065), .A1N(n1120), .B0(in_valid2), .Y(n1123) );
  AOI2BB2X1 U5550 ( .B0(in_valid), .B1(n5860), .A0N(n1038), .A1N(n873), .Y(
        n1124) );
  CLKINVX3 U5551 ( .A(in_valid2), .Y(n5833) );
  OAI22X1 U5552 ( .A0(n5074), .A1(n545), .B0(n5466), .B1(n4985), .Y(n4139) );
  OAI22X1 U5553 ( .A0(n5076), .A1(n513), .B0(n5488), .B1(n4985), .Y(n4011) );
  OAI22X1 U5554 ( .A0(n5077), .A1(n433), .B0(n5543), .B1(n4985), .Y(n3691) );
  OAI22X1 U5555 ( .A0(n5078), .A1(n385), .B0(n5578), .B1(n4985), .Y(n3563) );
  OAI22X1 U5556 ( .A0(n5074), .A1(n535), .B0(n5466), .B1(n4984), .Y(n4129) );
  OAI22X1 U5557 ( .A0(n5076), .A1(n503), .B0(n5488), .B1(n4984), .Y(n4001) );
  OAI22X1 U5558 ( .A0(n5077), .A1(n423), .B0(n5543), .B1(n4984), .Y(n3681) );
  OAI22X1 U5559 ( .A0(n5078), .A1(n375), .B0(n5578), .B1(n4984), .Y(n3553) );
  OAI22X1 U5560 ( .A0(n5074), .A1(n534), .B0(n5466), .B1(n4983), .Y(n4128) );
  OAI22X1 U5561 ( .A0(n5076), .A1(n502), .B0(n5488), .B1(n4983), .Y(n4000) );
  OAI22X1 U5562 ( .A0(n5077), .A1(n422), .B0(n5543), .B1(n4983), .Y(n3680) );
  OAI22X1 U5563 ( .A0(n5078), .A1(n374), .B0(n5578), .B1(n4983), .Y(n3552) );
  OAI22X1 U5564 ( .A0(n5074), .A1(n533), .B0(n5466), .B1(n4982), .Y(n4127) );
  OAI22X1 U5565 ( .A0(n5076), .A1(n501), .B0(n5488), .B1(n4982), .Y(n3999) );
  OAI22X1 U5566 ( .A0(n5077), .A1(n421), .B0(n5543), .B1(n4982), .Y(n3679) );
  OAI22X1 U5567 ( .A0(n5078), .A1(n373), .B0(n5578), .B1(n4982), .Y(n3551) );
  OAI22X1 U5568 ( .A0(n5074), .A1(n532), .B0(n5466), .B1(n4981), .Y(n4126) );
  OAI22X1 U5569 ( .A0(n5076), .A1(n500), .B0(n5488), .B1(n4981), .Y(n3998) );
  OAI22X1 U5570 ( .A0(n5077), .A1(n420), .B0(n5543), .B1(n4981), .Y(n3678) );
  OAI22X1 U5571 ( .A0(n5078), .A1(n372), .B0(n5578), .B1(n4981), .Y(n3550) );
  OAI22X1 U5572 ( .A0(n5074), .A1(n531), .B0(n5465), .B1(n4980), .Y(n4125) );
  OAI22X1 U5573 ( .A0(n5076), .A1(n499), .B0(n5487), .B1(n4980), .Y(n3997) );
  OAI22X1 U5574 ( .A0(n5077), .A1(n419), .B0(n5542), .B1(n4980), .Y(n3677) );
  OAI22X1 U5575 ( .A0(n5078), .A1(n371), .B0(n5577), .B1(n4980), .Y(n3549) );
  OAI22X1 U5576 ( .A0(n5074), .A1(n530), .B0(n5466), .B1(n4979), .Y(n4124) );
  OAI22X1 U5577 ( .A0(n5076), .A1(n498), .B0(n5488), .B1(n4979), .Y(n3996) );
  OAI22X1 U5578 ( .A0(n5077), .A1(n418), .B0(n5543), .B1(n4979), .Y(n3676) );
  OAI22X1 U5579 ( .A0(n5078), .A1(n370), .B0(n5578), .B1(n4979), .Y(n3548) );
  OAI22X1 U5580 ( .A0(n5336), .A1(n657), .B0(n5420), .B1(n4978), .Y(n4379) );
  OAI22X1 U5581 ( .A0(n5349), .A1(n609), .B0(n5442), .B1(n4978), .Y(n4251) );
  OAI22X1 U5582 ( .A0(n5377), .A1(n497), .B0(n5499), .B1(n4978), .Y(n3931) );
  OAI22X1 U5583 ( .A0(n5399), .A1(n465), .B0(n5521), .B1(n4978), .Y(n3803) );
  OAI22X1 U5584 ( .A0(n5336), .A1(n656), .B0(n5422), .B1(n4977), .Y(n4378) );
  OAI22X1 U5585 ( .A0(n5349), .A1(n608), .B0(n5444), .B1(n4977), .Y(n4250) );
  OAI22X1 U5586 ( .A0(n5377), .A1(n496), .B0(n5499), .B1(n4977), .Y(n3930) );
  OAI22X1 U5587 ( .A0(n5399), .A1(n464), .B0(n5521), .B1(n4977), .Y(n3802) );
  OAI22X1 U5588 ( .A0(n5336), .A1(n655), .B0(n5422), .B1(n4976), .Y(n4377) );
  OAI22X1 U5589 ( .A0(n5349), .A1(n607), .B0(n5444), .B1(n4976), .Y(n4249) );
  OAI22X1 U5590 ( .A0(n5376), .A1(n495), .B0(n5499), .B1(n4976), .Y(n3929) );
  OAI22X1 U5591 ( .A0(n5398), .A1(n463), .B0(n5521), .B1(n4976), .Y(n3801) );
  OAI22X1 U5592 ( .A0(n5336), .A1(n654), .B0(n5422), .B1(n4975), .Y(n4376) );
  OAI22X1 U5593 ( .A0(n5349), .A1(n606), .B0(n5444), .B1(n4975), .Y(n4248) );
  OAI22X1 U5594 ( .A0(n5376), .A1(n494), .B0(n5499), .B1(n4975), .Y(n3928) );
  OAI22X1 U5595 ( .A0(n5398), .A1(n462), .B0(n5521), .B1(n4975), .Y(n3800) );
  OAI22X1 U5596 ( .A0(n5074), .A1(n544), .B0(n5466), .B1(n4974), .Y(n4138) );
  OAI22X1 U5597 ( .A0(n5076), .A1(n512), .B0(n5488), .B1(n4974), .Y(n4010) );
  OAI22X1 U5598 ( .A0(n5077), .A1(n432), .B0(n5543), .B1(n4974), .Y(n3690) );
  OAI22X1 U5599 ( .A0(n5078), .A1(n384), .B0(n5578), .B1(n4974), .Y(n3562) );
  OAI22X1 U5600 ( .A0(n5336), .A1(n653), .B0(n5422), .B1(n4973), .Y(n4375) );
  OAI22X1 U5601 ( .A0(n5349), .A1(n605), .B0(n5444), .B1(n4973), .Y(n4247) );
  OAI22X1 U5602 ( .A0(n5369), .A1(n493), .B0(n5499), .B1(n4973), .Y(n3927) );
  OAI22X1 U5603 ( .A0(n5391), .A1(n461), .B0(n5521), .B1(n4973), .Y(n3799) );
  OAI22X1 U5604 ( .A0(n5336), .A1(n652), .B0(n5415), .B1(n4972), .Y(n4374) );
  OAI22X1 U5605 ( .A0(n5349), .A1(n604), .B0(n5437), .B1(n4972), .Y(n4246) );
  OAI22X1 U5606 ( .A0(n5370), .A1(n492), .B0(n5499), .B1(n4972), .Y(n3926) );
  OAI22X1 U5607 ( .A0(n5392), .A1(n460), .B0(n5521), .B1(n4972), .Y(n3798) );
  OAI22X1 U5608 ( .A0(n5336), .A1(n651), .B0(n5415), .B1(n4971), .Y(n4373) );
  OAI22X1 U5609 ( .A0(n5349), .A1(n603), .B0(n5437), .B1(n4971), .Y(n4245) );
  OAI22X1 U5610 ( .A0(n5375), .A1(n491), .B0(n5499), .B1(n4971), .Y(n3925) );
  OAI22X1 U5611 ( .A0(n5397), .A1(n459), .B0(n5521), .B1(n4971), .Y(n3797) );
  OAI22X1 U5612 ( .A0(n5336), .A1(n650), .B0(n5421), .B1(n4970), .Y(n4372) );
  OAI22X1 U5613 ( .A0(n5349), .A1(n602), .B0(n5443), .B1(n4970), .Y(n4244) );
  OAI22X1 U5614 ( .A0(n5375), .A1(n490), .B0(n5499), .B1(n4970), .Y(n3924) );
  OAI22X1 U5615 ( .A0(n5397), .A1(n458), .B0(n5521), .B1(n4970), .Y(n3796) );
  OAI22X1 U5616 ( .A0(n5336), .A1(n649), .B0(n5415), .B1(n4969), .Y(n4371) );
  OAI22X1 U5617 ( .A0(n5349), .A1(n601), .B0(n5437), .B1(n4969), .Y(n4243) );
  OAI22X1 U5618 ( .A0(n5374), .A1(n489), .B0(n5499), .B1(n4969), .Y(n3923) );
  OAI22X1 U5619 ( .A0(n5396), .A1(n457), .B0(n5521), .B1(n4969), .Y(n3795) );
  OAI22X1 U5620 ( .A0(n5336), .A1(n648), .B0(n5420), .B1(n4968), .Y(n4370) );
  OAI22X1 U5621 ( .A0(n5349), .A1(n600), .B0(n5442), .B1(n4968), .Y(n4242) );
  OAI22X1 U5622 ( .A0(n5374), .A1(n488), .B0(n5499), .B1(n4968), .Y(n3922) );
  OAI22X1 U5623 ( .A0(n5396), .A1(n456), .B0(n5521), .B1(n4968), .Y(n3794) );
  OAI22X1 U5624 ( .A0(n5336), .A1(n647), .B0(n5418), .B1(n4967), .Y(n4369) );
  OAI22X1 U5625 ( .A0(n5349), .A1(n599), .B0(n5440), .B1(n4967), .Y(n4241) );
  OAI22X1 U5626 ( .A0(n5373), .A1(n487), .B0(n5499), .B1(n4967), .Y(n3921) );
  OAI22X1 U5627 ( .A0(n5395), .A1(n455), .B0(n5521), .B1(n4967), .Y(n3793) );
  OAI22X1 U5628 ( .A0(n5336), .A1(n646), .B0(n5419), .B1(n4966), .Y(n4368) );
  OAI22X1 U5629 ( .A0(n5349), .A1(n598), .B0(n5441), .B1(n4966), .Y(n4240) );
  OAI22X1 U5630 ( .A0(n5373), .A1(n486), .B0(n5499), .B1(n4966), .Y(n3920) );
  OAI22X1 U5631 ( .A0(n5395), .A1(n454), .B0(n5521), .B1(n4966), .Y(n3792) );
  OAI22X1 U5632 ( .A0(n5335), .A1(n645), .B0(n5416), .B1(n4965), .Y(n4367) );
  OAI22X1 U5633 ( .A0(n5348), .A1(n597), .B0(n5438), .B1(n4965), .Y(n4239) );
  OAI22X1 U5634 ( .A0(n5377), .A1(n485), .B0(n5499), .B1(n4965), .Y(n3919) );
  OAI22X1 U5635 ( .A0(n5399), .A1(n453), .B0(n5521), .B1(n4965), .Y(n3791) );
  OAI22X1 U5636 ( .A0(n5335), .A1(n644), .B0(n5422), .B1(n4964), .Y(n4366) );
  OAI22X1 U5637 ( .A0(n5348), .A1(n596), .B0(n5444), .B1(n4964), .Y(n4238) );
  OAI22X1 U5638 ( .A0(n5373), .A1(n484), .B0(n5498), .B1(n4964), .Y(n3918) );
  OAI22X1 U5639 ( .A0(n5395), .A1(n452), .B0(n5520), .B1(n4964), .Y(n3790) );
  OAI22X1 U5640 ( .A0(n5074), .A1(n543), .B0(n5466), .B1(n4963), .Y(n4137) );
  OAI22X1 U5641 ( .A0(n5076), .A1(n511), .B0(n5488), .B1(n4963), .Y(n4009) );
  OAI22X1 U5642 ( .A0(n5077), .A1(n431), .B0(n5543), .B1(n4963), .Y(n3689) );
  OAI22X1 U5643 ( .A0(n5078), .A1(n383), .B0(n5578), .B1(n4963), .Y(n3561) );
  OAI22X1 U5644 ( .A0(n5335), .A1(n643), .B0(n5422), .B1(n4962), .Y(n4365) );
  OAI22X1 U5645 ( .A0(n5348), .A1(n595), .B0(n5444), .B1(n4962), .Y(n4237) );
  OAI22X1 U5646 ( .A0(n5372), .A1(n483), .B0(n5498), .B1(n4962), .Y(n3917) );
  OAI22X1 U5647 ( .A0(n5394), .A1(n451), .B0(n5520), .B1(n4962), .Y(n3789) );
  OAI22X1 U5648 ( .A0(n5335), .A1(n642), .B0(n5422), .B1(n4961), .Y(n4364) );
  OAI22X1 U5649 ( .A0(n5348), .A1(n594), .B0(n5444), .B1(n4961), .Y(n4236) );
  OAI22X1 U5650 ( .A0(n5372), .A1(n482), .B0(n5498), .B1(n4961), .Y(n3916) );
  OAI22X1 U5651 ( .A0(n5394), .A1(n450), .B0(n5520), .B1(n4961), .Y(n3788) );
  OAI22X1 U5652 ( .A0(n5074), .A1(n542), .B0(n5466), .B1(n4952), .Y(n4136) );
  OAI22X1 U5653 ( .A0(n5076), .A1(n510), .B0(n5488), .B1(n4952), .Y(n4008) );
  OAI22X1 U5654 ( .A0(n5077), .A1(n430), .B0(n5543), .B1(n4952), .Y(n3688) );
  OAI22X1 U5655 ( .A0(n5078), .A1(n382), .B0(n5578), .B1(n4952), .Y(n3560) );
  OAI22X1 U5656 ( .A0(n5074), .A1(n541), .B0(n5466), .B1(n4941), .Y(n4135) );
  OAI22X1 U5657 ( .A0(n5076), .A1(n509), .B0(n5488), .B1(n4941), .Y(n4007) );
  OAI22X1 U5658 ( .A0(n5077), .A1(n429), .B0(n5543), .B1(n4941), .Y(n3687) );
  OAI22X1 U5659 ( .A0(n5078), .A1(n381), .B0(n5578), .B1(n4941), .Y(n3559) );
  OAI22X1 U5660 ( .A0(n5074), .A1(n540), .B0(n5466), .B1(n4930), .Y(n4134) );
  OAI22X1 U5661 ( .A0(n5076), .A1(n508), .B0(n5488), .B1(n4930), .Y(n4006) );
  OAI22X1 U5662 ( .A0(n5077), .A1(n428), .B0(n5543), .B1(n4930), .Y(n3686) );
  OAI22X1 U5663 ( .A0(n5078), .A1(n380), .B0(n5578), .B1(n4930), .Y(n3558) );
  OAI22X1 U5664 ( .A0(n5074), .A1(n539), .B0(n5466), .B1(n4925), .Y(n4133) );
  OAI22X1 U5665 ( .A0(n5076), .A1(n507), .B0(n5488), .B1(n4925), .Y(n4005) );
  OAI22X1 U5666 ( .A0(n5077), .A1(n427), .B0(n5543), .B1(n4925), .Y(n3685) );
  OAI22X1 U5667 ( .A0(n5078), .A1(n379), .B0(n5578), .B1(n4925), .Y(n3557) );
  OAI22X1 U5668 ( .A0(n5074), .A1(n538), .B0(n5466), .B1(n4924), .Y(n4132) );
  OAI22X1 U5669 ( .A0(n5076), .A1(n506), .B0(n5488), .B1(n4924), .Y(n4004) );
  OAI22X1 U5670 ( .A0(n5077), .A1(n426), .B0(n5543), .B1(n4924), .Y(n3684) );
  OAI22X1 U5671 ( .A0(n5078), .A1(n378), .B0(n5578), .B1(n4924), .Y(n3556) );
  OAI22X1 U5672 ( .A0(n5074), .A1(n537), .B0(n5466), .B1(n4923), .Y(n4131) );
  OAI22X1 U5673 ( .A0(n5076), .A1(n505), .B0(n5488), .B1(n4923), .Y(n4003) );
  OAI22X1 U5674 ( .A0(n5077), .A1(n425), .B0(n5543), .B1(n4923), .Y(n3683) );
  OAI22X1 U5675 ( .A0(n5078), .A1(n377), .B0(n5578), .B1(n4923), .Y(n3555) );
  OAI22X1 U5676 ( .A0(n5074), .A1(n536), .B0(n5466), .B1(n4922), .Y(n4130) );
  OAI22X1 U5677 ( .A0(n5076), .A1(n504), .B0(n5488), .B1(n4922), .Y(n4002) );
  OAI22X1 U5678 ( .A0(n5077), .A1(n424), .B0(n5543), .B1(n4922), .Y(n3682) );
  OAI22X1 U5679 ( .A0(n5078), .A1(n376), .B0(n5578), .B1(n4922), .Y(n3554) );
  OAI22X1 U5680 ( .A0(n5073), .A1(n546), .B0(n5454), .B1(n4926), .Y(n4140) );
  OAI22X1 U5681 ( .A0(n5075), .A1(n514), .B0(n5476), .B1(n4926), .Y(n4012) );
  OAI22X1 U5682 ( .A0(n5369), .A1(n471), .B0(n5497), .B1(n4949), .Y(n3905) );
  OAI22X1 U5683 ( .A0(n5391), .A1(n439), .B0(n5519), .B1(n4949), .Y(n3777) );
  OAI22X1 U5684 ( .A0(n5369), .A1(n470), .B0(n5497), .B1(n4948), .Y(n3904) );
  OAI22X1 U5685 ( .A0(n5391), .A1(n438), .B0(n5519), .B1(n4948), .Y(n3776) );
  OAI22X1 U5686 ( .A0(n5368), .A1(n469), .B0(n5497), .B1(n4947), .Y(n3903) );
  OAI22X1 U5687 ( .A0(n5390), .A1(n437), .B0(n5519), .B1(n4947), .Y(n3775) );
  OAI22X1 U5688 ( .A0(n5368), .A1(n468), .B0(n5497), .B1(n4946), .Y(n3902) );
  OAI22X1 U5689 ( .A0(n5390), .A1(n436), .B0(n5519), .B1(n4946), .Y(n3774) );
  OAI22X1 U5690 ( .A0(n5369), .A1(n467), .B0(n5497), .B1(n4945), .Y(n3901) );
  OAI22X1 U5691 ( .A0(n5391), .A1(n435), .B0(n5519), .B1(n4945), .Y(n3773) );
  OAI22X1 U5692 ( .A0(n5368), .A1(n466), .B0(n5497), .B1(n4944), .Y(n3900) );
  OAI22X1 U5693 ( .A0(n5390), .A1(n434), .B0(n5519), .B1(n4944), .Y(n3772) );
  OAI22X1 U5694 ( .A0(n5335), .A1(n641), .B0(n5420), .B1(n4960), .Y(n4363) );
  OAI22X1 U5695 ( .A0(n5348), .A1(n593), .B0(n5442), .B1(n4960), .Y(n4235) );
  OAI22X1 U5696 ( .A0(n5370), .A1(n481), .B0(n5498), .B1(n4960), .Y(n3915) );
  OAI22X1 U5697 ( .A0(n5392), .A1(n449), .B0(n5520), .B1(n4960), .Y(n3787) );
  OAI22X1 U5698 ( .A0(n5335), .A1(n640), .B0(n5422), .B1(n4959), .Y(n4362) );
  OAI22X1 U5699 ( .A0(n5348), .A1(n592), .B0(n5444), .B1(n4959), .Y(n4234) );
  OAI22X1 U5700 ( .A0(n5376), .A1(n480), .B0(n5498), .B1(n4959), .Y(n3914) );
  OAI22X1 U5701 ( .A0(n5398), .A1(n448), .B0(n5520), .B1(n4959), .Y(n3786) );
  OAI22X1 U5702 ( .A0(n5335), .A1(n639), .B0(n5422), .B1(n4958), .Y(n4361) );
  OAI22X1 U5703 ( .A0(n5348), .A1(n591), .B0(n5444), .B1(n4958), .Y(n4233) );
  OAI22X1 U5704 ( .A0(n5377), .A1(n479), .B0(n5498), .B1(n4958), .Y(n3913) );
  OAI22X1 U5705 ( .A0(n5399), .A1(n447), .B0(n5520), .B1(n4958), .Y(n3785) );
  OAI22X1 U5706 ( .A0(n5335), .A1(n638), .B0(n5422), .B1(n4957), .Y(n4360) );
  OAI22X1 U5707 ( .A0(n5348), .A1(n590), .B0(n5444), .B1(n4957), .Y(n4232) );
  OAI22X1 U5708 ( .A0(n5373), .A1(n478), .B0(n5498), .B1(n4957), .Y(n3912) );
  OAI22X1 U5709 ( .A0(n5395), .A1(n446), .B0(n5520), .B1(n4957), .Y(n3784) );
  OAI22X1 U5710 ( .A0(n5335), .A1(n637), .B0(n5422), .B1(n4956), .Y(n4359) );
  OAI22X1 U5711 ( .A0(n5348), .A1(n589), .B0(n5444), .B1(n4956), .Y(n4231) );
  OAI22X1 U5712 ( .A0(n5371), .A1(n477), .B0(n5498), .B1(n4956), .Y(n3911) );
  OAI22X1 U5713 ( .A0(n5393), .A1(n445), .B0(n5520), .B1(n4956), .Y(n3783) );
  OAI22X1 U5714 ( .A0(n5335), .A1(n636), .B0(n5422), .B1(n4955), .Y(n4358) );
  OAI22X1 U5715 ( .A0(n5348), .A1(n588), .B0(n5444), .B1(n4955), .Y(n4230) );
  OAI22X1 U5716 ( .A0(n5371), .A1(n476), .B0(n5498), .B1(n4955), .Y(n3910) );
  OAI22X1 U5717 ( .A0(n5393), .A1(n444), .B0(n5520), .B1(n4955), .Y(n3782) );
  OAI22X1 U5718 ( .A0(n5335), .A1(n635), .B0(n5422), .B1(n4954), .Y(n4357) );
  OAI22X1 U5719 ( .A0(n5348), .A1(n587), .B0(n5444), .B1(n4954), .Y(n4229) );
  OAI22X1 U5720 ( .A0(n5370), .A1(n475), .B0(n5498), .B1(n4954), .Y(n3909) );
  OAI22X1 U5721 ( .A0(n5392), .A1(n443), .B0(n5520), .B1(n4954), .Y(n3781) );
  OAI22X1 U5722 ( .A0(n5335), .A1(n634), .B0(n5422), .B1(n4953), .Y(n4356) );
  OAI22X1 U5723 ( .A0(n5348), .A1(n586), .B0(n5444), .B1(n4953), .Y(n4228) );
  OAI22X1 U5724 ( .A0(n5370), .A1(n474), .B0(n5498), .B1(n4953), .Y(n3908) );
  OAI22X1 U5725 ( .A0(n5392), .A1(n442), .B0(n5520), .B1(n4953), .Y(n3780) );
  OAI22X1 U5726 ( .A0(n5334), .A1(n633), .B0(n5422), .B1(n4951), .Y(n4355) );
  OAI22X1 U5727 ( .A0(n5347), .A1(n585), .B0(n5444), .B1(n4951), .Y(n4227) );
  OAI22X1 U5728 ( .A0(n5375), .A1(n473), .B0(n5498), .B1(n4951), .Y(n3907) );
  OAI22X1 U5729 ( .A0(n5397), .A1(n441), .B0(n5520), .B1(n4951), .Y(n3779) );
  OAI22X1 U5730 ( .A0(n5334), .A1(n632), .B0(n5422), .B1(n4950), .Y(n4354) );
  OAI22X1 U5731 ( .A0(n5347), .A1(n584), .B0(n5444), .B1(n4950), .Y(n4226) );
  OAI22X1 U5732 ( .A0(n5374), .A1(n472), .B0(n5498), .B1(n4950), .Y(n3906) );
  OAI22X1 U5733 ( .A0(n5396), .A1(n440), .B0(n5520), .B1(n4950), .Y(n3778) );
  OAI22X1 U5734 ( .A0(n5334), .A1(n631), .B0(n5422), .B1(n4949), .Y(n4353) );
  OAI22X1 U5735 ( .A0(n5347), .A1(n583), .B0(n5444), .B1(n4949), .Y(n4225) );
  OAI22X1 U5736 ( .A0(n5334), .A1(n630), .B0(n5421), .B1(n4948), .Y(n4352) );
  OAI22X1 U5737 ( .A0(n5347), .A1(n582), .B0(n5443), .B1(n4948), .Y(n4224) );
  OAI22X1 U5738 ( .A0(n5334), .A1(n629), .B0(n5421), .B1(n4947), .Y(n4351) );
  OAI22X1 U5739 ( .A0(n5347), .A1(n581), .B0(n5443), .B1(n4947), .Y(n4223) );
  OAI22X1 U5740 ( .A0(n5334), .A1(n628), .B0(n5421), .B1(n4946), .Y(n4350) );
  OAI22X1 U5741 ( .A0(n5347), .A1(n580), .B0(n5443), .B1(n4946), .Y(n4222) );
  OAI22X1 U5742 ( .A0(n5334), .A1(n627), .B0(n5421), .B1(n4945), .Y(n4349) );
  OAI22X1 U5743 ( .A0(n5347), .A1(n579), .B0(n5443), .B1(n4945), .Y(n4221) );
  OAI22X1 U5744 ( .A0(n5334), .A1(n626), .B0(n5421), .B1(n4944), .Y(n4348) );
  OAI22X1 U5745 ( .A0(n5347), .A1(n578), .B0(n5443), .B1(n4944), .Y(n4220) );
  OAI22X1 U5746 ( .A0(n5334), .A1(n625), .B0(n5421), .B1(n4943), .Y(n4347) );
  OAI22X1 U5747 ( .A0(n5347), .A1(n577), .B0(n5443), .B1(n4943), .Y(n4219) );
  OAI22X1 U5748 ( .A0(n5073), .A1(n561), .B0(n5455), .B1(n4943), .Y(n4155) );
  OAI22X1 U5749 ( .A0(n5075), .A1(n529), .B0(n5477), .B1(n4943), .Y(n4027) );
  OAI22X1 U5750 ( .A0(n5334), .A1(n624), .B0(n5421), .B1(n4942), .Y(n4346) );
  OAI22X1 U5751 ( .A0(n5347), .A1(n576), .B0(n5443), .B1(n4942), .Y(n4218) );
  OAI22X1 U5752 ( .A0(n5073), .A1(n560), .B0(n5455), .B1(n4942), .Y(n4154) );
  OAI22X1 U5753 ( .A0(n5075), .A1(n528), .B0(n5477), .B1(n4942), .Y(n4026) );
  OAI22X1 U5754 ( .A0(n5334), .A1(n623), .B0(n5421), .B1(n4940), .Y(n4345) );
  OAI22X1 U5755 ( .A0(n5347), .A1(n575), .B0(n5443), .B1(n4940), .Y(n4217) );
  OAI22X1 U5756 ( .A0(n5073), .A1(n559), .B0(n5455), .B1(n4940), .Y(n4153) );
  OAI22X1 U5757 ( .A0(n5075), .A1(n527), .B0(n5477), .B1(n4940), .Y(n4025) );
  OAI22X1 U5758 ( .A0(n5334), .A1(n622), .B0(n5421), .B1(n4939), .Y(n4344) );
  OAI22X1 U5759 ( .A0(n5347), .A1(n574), .B0(n5443), .B1(n4939), .Y(n4216) );
  OAI22X1 U5760 ( .A0(n5073), .A1(n558), .B0(n5455), .B1(n4939), .Y(n4152) );
  OAI22X1 U5761 ( .A0(n5075), .A1(n526), .B0(n5477), .B1(n4939), .Y(n4024) );
  OAI22X1 U5762 ( .A0(n5334), .A1(n621), .B0(n5421), .B1(n4938), .Y(n4343) );
  OAI22X1 U5763 ( .A0(n5347), .A1(n573), .B0(n5443), .B1(n4938), .Y(n4215) );
  OAI22X1 U5764 ( .A0(n5073), .A1(n557), .B0(n5455), .B1(n4938), .Y(n4151) );
  OAI22X1 U5765 ( .A0(n5075), .A1(n525), .B0(n5477), .B1(n4938), .Y(n4023) );
  OAI22X1 U5766 ( .A0(n5334), .A1(n620), .B0(n5421), .B1(n4937), .Y(n4342) );
  OAI22X1 U5767 ( .A0(n5347), .A1(n572), .B0(n5443), .B1(n4937), .Y(n4214) );
  OAI22X1 U5768 ( .A0(n5073), .A1(n556), .B0(n5455), .B1(n4937), .Y(n4150) );
  OAI22X1 U5769 ( .A0(n5075), .A1(n524), .B0(n5477), .B1(n4937), .Y(n4022) );
  OAI22X1 U5770 ( .A0(n5334), .A1(n619), .B0(n5421), .B1(n4936), .Y(n4341) );
  OAI22X1 U5771 ( .A0(n5347), .A1(n571), .B0(n5443), .B1(n4936), .Y(n4213) );
  OAI22X1 U5772 ( .A0(n5073), .A1(n555), .B0(n5455), .B1(n4936), .Y(n4149) );
  OAI22X1 U5773 ( .A0(n5075), .A1(n523), .B0(n5477), .B1(n4936), .Y(n4021) );
  OAI22X1 U5774 ( .A0(n5334), .A1(n618), .B0(n5421), .B1(n4935), .Y(n4340) );
  OAI22X1 U5775 ( .A0(n5347), .A1(n570), .B0(n5443), .B1(n4935), .Y(n4212) );
  OAI22X1 U5776 ( .A0(n5073), .A1(n554), .B0(n5455), .B1(n4935), .Y(n4148) );
  OAI22X1 U5777 ( .A0(n5075), .A1(n522), .B0(n5477), .B1(n4935), .Y(n4020) );
  OAI22X1 U5778 ( .A0(n5334), .A1(n617), .B0(n5420), .B1(n4934), .Y(n4339) );
  OAI22X1 U5779 ( .A0(n5347), .A1(n569), .B0(n5442), .B1(n4934), .Y(n4211) );
  OAI22X1 U5780 ( .A0(n5073), .A1(n553), .B0(n5455), .B1(n4934), .Y(n4147) );
  OAI22X1 U5781 ( .A0(n5075), .A1(n521), .B0(n5477), .B1(n4934), .Y(n4019) );
  OAI22X1 U5782 ( .A0(n5336), .A1(n616), .B0(n5420), .B1(n4933), .Y(n4338) );
  OAI22X1 U5783 ( .A0(n5349), .A1(n568), .B0(n5442), .B1(n4933), .Y(n4210) );
  OAI22X1 U5784 ( .A0(n5073), .A1(n552), .B0(n5455), .B1(n4933), .Y(n4146) );
  OAI22X1 U5785 ( .A0(n5075), .A1(n520), .B0(n5477), .B1(n4933), .Y(n4018) );
  OAI22X1 U5786 ( .A0(n5335), .A1(n615), .B0(n5420), .B1(n4932), .Y(n4337) );
  OAI22X1 U5787 ( .A0(n5348), .A1(n567), .B0(n5442), .B1(n4932), .Y(n4209) );
  OAI22X1 U5788 ( .A0(n5073), .A1(n551), .B0(n5455), .B1(n4932), .Y(n4145) );
  OAI22X1 U5789 ( .A0(n5075), .A1(n519), .B0(n5477), .B1(n4932), .Y(n4017) );
  OAI22X1 U5790 ( .A0(n5336), .A1(n614), .B0(n5420), .B1(n4931), .Y(n4336) );
  OAI22X1 U5791 ( .A0(n5349), .A1(n566), .B0(n5442), .B1(n4931), .Y(n4208) );
  OAI22X1 U5792 ( .A0(n5073), .A1(n550), .B0(n5455), .B1(n4931), .Y(n4144) );
  OAI22X1 U5793 ( .A0(n5075), .A1(n518), .B0(n5477), .B1(n4931), .Y(n4016) );
  OAI22X1 U5794 ( .A0(n5335), .A1(n613), .B0(n5420), .B1(n4929), .Y(n4335) );
  OAI22X1 U5795 ( .A0(n5348), .A1(n565), .B0(n5442), .B1(n4929), .Y(n4207) );
  OAI22X1 U5796 ( .A0(n5073), .A1(n549), .B0(n5455), .B1(n4929), .Y(n4143) );
  OAI22X1 U5797 ( .A0(n5075), .A1(n517), .B0(n5477), .B1(n4929), .Y(n4015) );
  OAI22X1 U5798 ( .A0(n5336), .A1(n612), .B0(n5420), .B1(n4928), .Y(n4334) );
  OAI22X1 U5799 ( .A0(n5349), .A1(n564), .B0(n5442), .B1(n4928), .Y(n4206) );
  OAI22X1 U5800 ( .A0(n5073), .A1(n548), .B0(n5455), .B1(n4928), .Y(n4142) );
  OAI22X1 U5801 ( .A0(n5075), .A1(n516), .B0(n5477), .B1(n4928), .Y(n4014) );
  OAI22X1 U5802 ( .A0(n5335), .A1(n611), .B0(n5420), .B1(n4927), .Y(n4333) );
  OAI22X1 U5803 ( .A0(n5348), .A1(n563), .B0(n5442), .B1(n4927), .Y(n4205) );
  OAI22X1 U5804 ( .A0(n5073), .A1(n547), .B0(n5455), .B1(n4927), .Y(n4141) );
  OAI22X1 U5805 ( .A0(n5075), .A1(n515), .B0(n5477), .B1(n4927), .Y(n4013) );
  OAI22X1 U5806 ( .A0(n5336), .A1(n610), .B0(n5420), .B1(n4926), .Y(n4332) );
  OAI22X1 U5807 ( .A0(n5349), .A1(n562), .B0(n5442), .B1(n4926), .Y(n4204) );
  AOI211X1 U5808 ( .A0(n1115), .A1(n5833), .B0(n1116), .C0(n5250), .Y(n1114)
         );
  AND4X2 U5809 ( .A(cs[2]), .B(n5858), .C(cs[1]), .D(cs[0]), .Y(n1116) );
  NAND3X1 U5810 ( .A(n5889), .B(n5858), .C(n1119), .Y(n1117) );
  OAI21XL U5811 ( .A0(in_valid), .A1(n5833), .B0(n5883), .Y(n1119) );
  OAI2BB2X1 U5812 ( .B0(n4992), .B1(n5405), .A0N(w_matrix[61]), .A1N(n5097), 
        .Y(n3374) );
  OAI2BB2X1 U5813 ( .B0(n4992), .B1(n5427), .A0N(w_matrix[189]), .A1N(n5107), 
        .Y(n3246) );
  OAI2BB2X1 U5814 ( .B0(n4992), .B1(n5504), .A0N(w_matrix[637]), .A1N(n5149), 
        .Y(n2798) );
  OAI2BB2X1 U5815 ( .B0(n4992), .B1(n5530), .A0N(w_matrix[765]), .A1N(n5151), 
        .Y(n2670) );
  OAI2BB2X1 U5816 ( .B0(n4991), .B1(n5406), .A0N(w_matrix[62]), .A1N(n5097), 
        .Y(n3373) );
  OAI2BB2X1 U5817 ( .B0(n4991), .B1(n5428), .A0N(w_matrix[190]), .A1N(n5107), 
        .Y(n3245) );
  OAI2BB2X1 U5818 ( .B0(n4991), .B1(n5505), .A0N(w_matrix[638]), .A1N(n5149), 
        .Y(n2797) );
  OAI2BB2X1 U5819 ( .B0(n4991), .B1(n5531), .A0N(w_matrix[766]), .A1N(n5151), 
        .Y(n2669) );
  OAI2BB2X1 U5820 ( .B0(n4990), .B1(n5404), .A0N(w_matrix[63]), .A1N(n5097), 
        .Y(n3372) );
  OAI2BB2X1 U5821 ( .B0(n4990), .B1(n5426), .A0N(w_matrix[191]), .A1N(n5107), 
        .Y(n3244) );
  OAI2BB2X1 U5822 ( .B0(n4990), .B1(n5503), .A0N(w_matrix[639]), .A1N(n5149), 
        .Y(n2796) );
  OAI2BB2X1 U5823 ( .B0(n4990), .B1(n5531), .A0N(w_matrix[767]), .A1N(n5151), 
        .Y(n2668) );
  OAI2BB2X1 U5824 ( .B0(n5408), .B1(n4985), .A0N(n5097), .A1N(x_matrix[0]), 
        .Y(n4459) );
  OAI2BB2X1 U5825 ( .B0(n5415), .B1(n4985), .A0N(n5338), .A1N(x_matrix[64]), 
        .Y(n4395) );
  OAI2BB2X1 U5826 ( .B0(n5430), .B1(n4985), .A0N(n5107), .A1N(x_matrix[80]), 
        .Y(n4331) );
  OAI2BB2X1 U5827 ( .B0(n5437), .B1(n4985), .A0N(n5351), .A1N(x_matrix[144]), 
        .Y(n4267) );
  OAI2BB2X1 U5828 ( .B0(n5448), .B1(n4985), .A0N(n5109), .A1N(x_matrix[160]), 
        .Y(n4203) );
  OAI2BB2X1 U5829 ( .B0(n5470), .B1(n4985), .A0N(n5125), .A1N(x_matrix[256]), 
        .Y(n4075) );
  OAI2BB2X1 U5830 ( .B0(n5492), .B1(n4985), .A0N(n5360), .A1N(x_matrix[352]), 
        .Y(n3947) );
  OAI2BB2X1 U5831 ( .B0(n5507), .B1(n4985), .A0N(n5149), .A1N(x_matrix[384]), 
        .Y(n3883) );
  OAI2BB2X1 U5832 ( .B0(n5514), .B1(n4985), .A0N(n5382), .A1N(x_matrix[448]), 
        .Y(n3819) );
  OAI2BB2X1 U5833 ( .B0(n5529), .B1(n4985), .A0N(n5151), .A1N(x_matrix[480]), 
        .Y(n3755) );
  OAI2BB2X1 U5834 ( .B0(n5411), .B1(n4984), .A0N(n5097), .A1N(x_matrix[10]), 
        .Y(n4449) );
  OAI2BB2X1 U5835 ( .B0(n5415), .B1(n4984), .A0N(n5341), .A1N(x_matrix[74]), 
        .Y(n4385) );
  OAI2BB2X1 U5836 ( .B0(n5433), .B1(n4984), .A0N(n5107), .A1N(x_matrix[90]), 
        .Y(n4321) );
  OAI2BB2X1 U5837 ( .B0(n5437), .B1(n4984), .A0N(n5354), .A1N(x_matrix[154]), 
        .Y(n4257) );
  OAI2BB2X1 U5838 ( .B0(n5448), .B1(n4984), .A0N(n5109), .A1N(x_matrix[170]), 
        .Y(n4193) );
  OAI2BB2X1 U5839 ( .B0(n5470), .B1(n4984), .A0N(n5125), .A1N(x_matrix[266]), 
        .Y(n4065) );
  OAI2BB2X1 U5840 ( .B0(n5492), .B1(n4984), .A0N(n5360), .A1N(x_matrix[362]), 
        .Y(n3937) );
  OAI2BB2X1 U5841 ( .B0(n5510), .B1(n4984), .A0N(n5149), .A1N(x_matrix[394]), 
        .Y(n3873) );
  OAI2BB2X1 U5842 ( .B0(n5514), .B1(n4984), .A0N(n5382), .A1N(x_matrix[458]), 
        .Y(n3809) );
  OAI2BB2X1 U5843 ( .B0(n5532), .B1(n4984), .A0N(n5151), .A1N(x_matrix[490]), 
        .Y(n3745) );
  OAI2BB2X1 U5844 ( .B0(n5408), .B1(n4983), .A0N(n5097), .A1N(x_matrix[11]), 
        .Y(n4448) );
  OAI2BB2X1 U5845 ( .B0(n5415), .B1(n4983), .A0N(n5344), .A1N(x_matrix[75]), 
        .Y(n4384) );
  OAI2BB2X1 U5846 ( .B0(n5430), .B1(n4983), .A0N(n5107), .A1N(x_matrix[91]), 
        .Y(n4320) );
  OAI2BB2X1 U5847 ( .B0(n5437), .B1(n4983), .A0N(n5357), .A1N(x_matrix[155]), 
        .Y(n4256) );
  OAI2BB2X1 U5848 ( .B0(n5448), .B1(n4983), .A0N(n5109), .A1N(x_matrix[171]), 
        .Y(n4192) );
  OAI2BB2X1 U5849 ( .B0(n5470), .B1(n4983), .A0N(n5125), .A1N(x_matrix[267]), 
        .Y(n4064) );
  OAI2BB2X1 U5850 ( .B0(n5492), .B1(n4983), .A0N(n5360), .A1N(x_matrix[363]), 
        .Y(n3936) );
  OAI2BB2X1 U5851 ( .B0(n5507), .B1(n4983), .A0N(n5149), .A1N(x_matrix[395]), 
        .Y(n3872) );
  OAI2BB2X1 U5852 ( .B0(n5514), .B1(n4983), .A0N(n5382), .A1N(x_matrix[459]), 
        .Y(n3808) );
  OAI2BB2X1 U5853 ( .B0(n5527), .B1(n4983), .A0N(n5151), .A1N(x_matrix[491]), 
        .Y(n3744) );
  OAI2BB2X1 U5854 ( .B0(n5404), .B1(n4982), .A0N(n5089), .A1N(x_matrix[12]), 
        .Y(n4447) );
  OAI2BB2X1 U5855 ( .B0(n5416), .B1(n4982), .A0N(n5341), .A1N(x_matrix[76]), 
        .Y(n4383) );
  OAI2BB2X1 U5856 ( .B0(n5426), .B1(n4982), .A0N(n5099), .A1N(x_matrix[92]), 
        .Y(n4319) );
  OAI2BB2X1 U5857 ( .B0(n5438), .B1(n4982), .A0N(n5354), .A1N(x_matrix[156]), 
        .Y(n4255) );
  OAI2BB2X1 U5858 ( .B0(n5449), .B1(n4982), .A0N(n5110), .A1N(x_matrix[172]), 
        .Y(n4191) );
  OAI2BB2X1 U5859 ( .B0(n5471), .B1(n4982), .A0N(n5126), .A1N(x_matrix[268]), 
        .Y(n4063) );
  OAI2BB2X1 U5860 ( .B0(n5492), .B1(n4982), .A0N(n5361), .A1N(x_matrix[364]), 
        .Y(n3935) );
  OAI2BB2X1 U5861 ( .B0(n5503), .B1(n4982), .A0N(n5141), .A1N(x_matrix[396]), 
        .Y(n3871) );
  OAI2BB2X1 U5862 ( .B0(n5514), .B1(n4982), .A0N(n5383), .A1N(x_matrix[460]), 
        .Y(n3807) );
  OAI2BB2X1 U5863 ( .B0(n5525), .B1(n4982), .A0N(n5152), .A1N(x_matrix[492]), 
        .Y(n3743) );
  OAI2BB2X1 U5864 ( .B0(n5404), .B1(n4981), .A0N(n5089), .A1N(x_matrix[13]), 
        .Y(n4446) );
  OAI2BB2X1 U5865 ( .B0(n5416), .B1(n4981), .A0N(n5343), .A1N(x_matrix[77]), 
        .Y(n4382) );
  OAI2BB2X1 U5866 ( .B0(n5426), .B1(n4981), .A0N(n5099), .A1N(x_matrix[93]), 
        .Y(n4318) );
  OAI2BB2X1 U5867 ( .B0(n5438), .B1(n4981), .A0N(n5356), .A1N(x_matrix[157]), 
        .Y(n4254) );
  OAI2BB2X1 U5868 ( .B0(n5449), .B1(n4981), .A0N(n5110), .A1N(x_matrix[173]), 
        .Y(n4190) );
  OAI2BB2X1 U5869 ( .B0(n5471), .B1(n4981), .A0N(n5126), .A1N(x_matrix[269]), 
        .Y(n4062) );
  OAI2BB2X1 U5870 ( .B0(n5499), .B1(n4981), .A0N(n5361), .A1N(x_matrix[365]), 
        .Y(n3934) );
  OAI2BB2X1 U5871 ( .B0(n5503), .B1(n4981), .A0N(n5141), .A1N(x_matrix[397]), 
        .Y(n3870) );
  OAI2BB2X1 U5872 ( .B0(n5521), .B1(n4981), .A0N(n5383), .A1N(x_matrix[461]), 
        .Y(n3806) );
  OAI2BB2X1 U5873 ( .B0(n5525), .B1(n4981), .A0N(n5152), .A1N(x_matrix[493]), 
        .Y(n3742) );
  OAI2BB2X1 U5874 ( .B0(n5404), .B1(n4980), .A0N(n5089), .A1N(x_matrix[14]), 
        .Y(n4445) );
  OAI2BB2X1 U5875 ( .B0(n5416), .B1(n4980), .A0N(n5341), .A1N(x_matrix[78]), 
        .Y(n4381) );
  OAI2BB2X1 U5876 ( .B0(n5426), .B1(n4980), .A0N(n5099), .A1N(x_matrix[94]), 
        .Y(n4317) );
  OAI2BB2X1 U5877 ( .B0(n5438), .B1(n4980), .A0N(n5354), .A1N(x_matrix[158]), 
        .Y(n4253) );
  OAI2BB2X1 U5878 ( .B0(n5449), .B1(n4980), .A0N(n5110), .A1N(x_matrix[174]), 
        .Y(n4189) );
  OAI2BB2X1 U5879 ( .B0(n5471), .B1(n4980), .A0N(n5126), .A1N(x_matrix[270]), 
        .Y(n4061) );
  OAI2BB2X1 U5880 ( .B0(n5498), .B1(n4980), .A0N(n5361), .A1N(x_matrix[366]), 
        .Y(n3933) );
  OAI2BB2X1 U5881 ( .B0(n5503), .B1(n4980), .A0N(n5141), .A1N(x_matrix[398]), 
        .Y(n3869) );
  OAI2BB2X1 U5882 ( .B0(n5520), .B1(n4980), .A0N(n5383), .A1N(x_matrix[462]), 
        .Y(n3805) );
  OAI2BB2X1 U5883 ( .B0(n5525), .B1(n4980), .A0N(n5152), .A1N(x_matrix[494]), 
        .Y(n3741) );
  OAI2BB2X1 U5884 ( .B0(n5404), .B1(n4979), .A0N(n5089), .A1N(x_matrix[15]), 
        .Y(n4444) );
  OAI2BB2X1 U5885 ( .B0(n5416), .B1(n4979), .A0N(n5344), .A1N(x_matrix[79]), 
        .Y(n4380) );
  OAI2BB2X1 U5886 ( .B0(n5426), .B1(n4979), .A0N(n5099), .A1N(x_matrix[95]), 
        .Y(n4316) );
  OAI2BB2X1 U5887 ( .B0(n5438), .B1(n4979), .A0N(n5357), .A1N(x_matrix[159]), 
        .Y(n4252) );
  OAI2BB2X1 U5888 ( .B0(n5449), .B1(n4979), .A0N(n5110), .A1N(x_matrix[175]), 
        .Y(n4188) );
  OAI2BB2X1 U5889 ( .B0(n5471), .B1(n4979), .A0N(n5126), .A1N(x_matrix[271]), 
        .Y(n4060) );
  OAI2BB2X1 U5890 ( .B0(n5492), .B1(n4979), .A0N(n5361), .A1N(x_matrix[367]), 
        .Y(n3932) );
  OAI2BB2X1 U5891 ( .B0(n5503), .B1(n4979), .A0N(n5141), .A1N(x_matrix[399]), 
        .Y(n3868) );
  OAI2BB2X1 U5892 ( .B0(n5514), .B1(n4979), .A0N(n5383), .A1N(x_matrix[463]), 
        .Y(n3804) );
  OAI2BB2X1 U5893 ( .B0(n5525), .B1(n4979), .A0N(n5152), .A1N(x_matrix[495]), 
        .Y(n3740) );
  OAI2BB2X1 U5894 ( .B0(n5411), .B1(n4974), .A0N(n5097), .A1N(x_matrix[1]), 
        .Y(n4458) );
  OAI2BB2X1 U5895 ( .B0(n5415), .B1(n4974), .A0N(n5337), .A1N(x_matrix[65]), 
        .Y(n4394) );
  OAI2BB2X1 U5896 ( .B0(n5433), .B1(n4974), .A0N(n5107), .A1N(x_matrix[81]), 
        .Y(n4330) );
  OAI2BB2X1 U5897 ( .B0(n5437), .B1(n4974), .A0N(n5350), .A1N(x_matrix[145]), 
        .Y(n4266) );
  OAI2BB2X1 U5898 ( .B0(n5448), .B1(n4974), .A0N(n5109), .A1N(x_matrix[161]), 
        .Y(n4202) );
  OAI2BB2X1 U5899 ( .B0(n5470), .B1(n4974), .A0N(n5125), .A1N(x_matrix[257]), 
        .Y(n4074) );
  OAI2BB2X1 U5900 ( .B0(n5492), .B1(n4974), .A0N(n5360), .A1N(x_matrix[353]), 
        .Y(n3946) );
  OAI2BB2X1 U5901 ( .B0(n5510), .B1(n4974), .A0N(n5149), .A1N(x_matrix[385]), 
        .Y(n3882) );
  OAI2BB2X1 U5902 ( .B0(n5514), .B1(n4974), .A0N(n5382), .A1N(x_matrix[449]), 
        .Y(n3818) );
  OAI2BB2X1 U5903 ( .B0(n5528), .B1(n4974), .A0N(n5151), .A1N(x_matrix[481]), 
        .Y(n3754) );
  OAI2BB2X1 U5904 ( .B0(n5408), .B1(n4963), .A0N(n5097), .A1N(x_matrix[2]), 
        .Y(n4457) );
  OAI2BB2X1 U5905 ( .B0(n5415), .B1(n4963), .A0N(n5344), .A1N(x_matrix[66]), 
        .Y(n4393) );
  OAI2BB2X1 U5906 ( .B0(n5430), .B1(n4963), .A0N(n5107), .A1N(x_matrix[82]), 
        .Y(n4329) );
  OAI2BB2X1 U5907 ( .B0(n5437), .B1(n4963), .A0N(n5357), .A1N(x_matrix[146]), 
        .Y(n4265) );
  OAI2BB2X1 U5908 ( .B0(n5448), .B1(n4963), .A0N(n5109), .A1N(x_matrix[162]), 
        .Y(n4201) );
  OAI2BB2X1 U5909 ( .B0(n5470), .B1(n4963), .A0N(n5125), .A1N(x_matrix[258]), 
        .Y(n4073) );
  OAI2BB2X1 U5910 ( .B0(n5492), .B1(n4963), .A0N(n5360), .A1N(x_matrix[354]), 
        .Y(n3945) );
  OAI2BB2X1 U5911 ( .B0(n5507), .B1(n4963), .A0N(n5149), .A1N(x_matrix[386]), 
        .Y(n3881) );
  OAI2BB2X1 U5912 ( .B0(n5514), .B1(n4963), .A0N(n5382), .A1N(x_matrix[450]), 
        .Y(n3817) );
  OAI2BB2X1 U5913 ( .B0(n5525), .B1(n4963), .A0N(n5151), .A1N(x_matrix[482]), 
        .Y(n3753) );
  OAI2BB2X1 U5914 ( .B0(n5411), .B1(n4952), .A0N(n5097), .A1N(x_matrix[3]), 
        .Y(n4456) );
  OAI2BB2X1 U5915 ( .B0(n5415), .B1(n4952), .A0N(n5338), .A1N(x_matrix[67]), 
        .Y(n4392) );
  OAI2BB2X1 U5916 ( .B0(n5433), .B1(n4952), .A0N(n5107), .A1N(x_matrix[83]), 
        .Y(n4328) );
  OAI2BB2X1 U5917 ( .B0(n5437), .B1(n4952), .A0N(n5351), .A1N(x_matrix[147]), 
        .Y(n4264) );
  OAI2BB2X1 U5918 ( .B0(n5448), .B1(n4952), .A0N(n5109), .A1N(x_matrix[163]), 
        .Y(n4200) );
  OAI2BB2X1 U5919 ( .B0(n5470), .B1(n4952), .A0N(n5125), .A1N(x_matrix[259]), 
        .Y(n4072) );
  OAI2BB2X1 U5920 ( .B0(n5492), .B1(n4952), .A0N(n5360), .A1N(x_matrix[355]), 
        .Y(n3944) );
  OAI2BB2X1 U5921 ( .B0(n5510), .B1(n4952), .A0N(n5149), .A1N(x_matrix[387]), 
        .Y(n3880) );
  OAI2BB2X1 U5922 ( .B0(n5514), .B1(n4952), .A0N(n5382), .A1N(x_matrix[451]), 
        .Y(n3816) );
  OAI2BB2X1 U5923 ( .B0(n5526), .B1(n4952), .A0N(n5151), .A1N(x_matrix[483]), 
        .Y(n3752) );
  OAI2BB2X1 U5924 ( .B0(n5408), .B1(n4941), .A0N(n5097), .A1N(x_matrix[4]), 
        .Y(n4455) );
  OAI2BB2X1 U5925 ( .B0(n5415), .B1(n4941), .A0N(n5342), .A1N(x_matrix[68]), 
        .Y(n4391) );
  OAI2BB2X1 U5926 ( .B0(n5430), .B1(n4941), .A0N(n5107), .A1N(x_matrix[84]), 
        .Y(n4327) );
  OAI2BB2X1 U5927 ( .B0(n5437), .B1(n4941), .A0N(n5355), .A1N(x_matrix[148]), 
        .Y(n4263) );
  OAI2BB2X1 U5928 ( .B0(n5448), .B1(n4941), .A0N(n5109), .A1N(x_matrix[164]), 
        .Y(n4199) );
  OAI2BB2X1 U5929 ( .B0(n5470), .B1(n4941), .A0N(n5125), .A1N(x_matrix[260]), 
        .Y(n4071) );
  OAI2BB2X1 U5930 ( .B0(n5492), .B1(n4941), .A0N(n5360), .A1N(x_matrix[356]), 
        .Y(n3943) );
  OAI2BB2X1 U5931 ( .B0(n5507), .B1(n4941), .A0N(n5149), .A1N(x_matrix[388]), 
        .Y(n3879) );
  OAI2BB2X1 U5932 ( .B0(n5514), .B1(n4941), .A0N(n5382), .A1N(x_matrix[452]), 
        .Y(n3815) );
  OAI2BB2X1 U5933 ( .B0(n5532), .B1(n4941), .A0N(n5151), .A1N(x_matrix[484]), 
        .Y(n3751) );
  OAI2BB2X1 U5934 ( .B0(n5411), .B1(n4930), .A0N(n5097), .A1N(x_matrix[5]), 
        .Y(n4454) );
  OAI2BB2X1 U5935 ( .B0(n5415), .B1(n4930), .A0N(n5343), .A1N(x_matrix[69]), 
        .Y(n4390) );
  OAI2BB2X1 U5936 ( .B0(n5433), .B1(n4930), .A0N(n5107), .A1N(x_matrix[85]), 
        .Y(n4326) );
  OAI2BB2X1 U5937 ( .B0(n5437), .B1(n4930), .A0N(n5356), .A1N(x_matrix[149]), 
        .Y(n4262) );
  OAI2BB2X1 U5938 ( .B0(n5448), .B1(n4930), .A0N(n5109), .A1N(x_matrix[165]), 
        .Y(n4198) );
  OAI2BB2X1 U5939 ( .B0(n5470), .B1(n4930), .A0N(n5125), .A1N(x_matrix[261]), 
        .Y(n4070) );
  OAI2BB2X1 U5940 ( .B0(n5492), .B1(n4930), .A0N(n5360), .A1N(x_matrix[357]), 
        .Y(n3942) );
  OAI2BB2X1 U5941 ( .B0(n5510), .B1(n4930), .A0N(n5149), .A1N(x_matrix[389]), 
        .Y(n3878) );
  OAI2BB2X1 U5942 ( .B0(n5514), .B1(n4930), .A0N(n5382), .A1N(x_matrix[453]), 
        .Y(n3814) );
  OAI2BB2X1 U5943 ( .B0(n5527), .B1(n4930), .A0N(n5151), .A1N(x_matrix[485]), 
        .Y(n3750) );
  OAI2BB2X1 U5944 ( .B0(n5409), .B1(n4925), .A0N(n5097), .A1N(x_matrix[6]), 
        .Y(n4453) );
  OAI2BB2X1 U5945 ( .B0(n5415), .B1(n4925), .A0N(n5343), .A1N(x_matrix[70]), 
        .Y(n4389) );
  OAI2BB2X1 U5946 ( .B0(n5431), .B1(n4925), .A0N(n5107), .A1N(x_matrix[86]), 
        .Y(n4325) );
  OAI2BB2X1 U5947 ( .B0(n5437), .B1(n4925), .A0N(n5356), .A1N(x_matrix[150]), 
        .Y(n4261) );
  OAI2BB2X1 U5948 ( .B0(n5448), .B1(n4925), .A0N(n5109), .A1N(x_matrix[166]), 
        .Y(n4197) );
  OAI2BB2X1 U5949 ( .B0(n5470), .B1(n4925), .A0N(n5125), .A1N(x_matrix[262]), 
        .Y(n4069) );
  OAI2BB2X1 U5950 ( .B0(n5492), .B1(n4925), .A0N(n5360), .A1N(x_matrix[358]), 
        .Y(n3941) );
  OAI2BB2X1 U5951 ( .B0(n5508), .B1(n4925), .A0N(n5149), .A1N(x_matrix[390]), 
        .Y(n3877) );
  OAI2BB2X1 U5952 ( .B0(n5514), .B1(n4925), .A0N(n5382), .A1N(x_matrix[454]), 
        .Y(n3813) );
  OAI2BB2X1 U5953 ( .B0(n5528), .B1(n4925), .A0N(n5151), .A1N(x_matrix[486]), 
        .Y(n3749) );
  OAI2BB2X1 U5954 ( .B0(n5410), .B1(n4924), .A0N(n5089), .A1N(x_matrix[7]), 
        .Y(n4452) );
  OAI2BB2X1 U5955 ( .B0(n5415), .B1(n4924), .A0N(n5343), .A1N(x_matrix[71]), 
        .Y(n4388) );
  OAI2BB2X1 U5956 ( .B0(n5432), .B1(n4924), .A0N(n5099), .A1N(x_matrix[87]), 
        .Y(n4324) );
  OAI2BB2X1 U5957 ( .B0(n5437), .B1(n4924), .A0N(n5356), .A1N(x_matrix[151]), 
        .Y(n4260) );
  OAI2BB2X1 U5958 ( .B0(n5448), .B1(n4924), .A0N(n5109), .A1N(x_matrix[167]), 
        .Y(n4196) );
  OAI2BB2X1 U5959 ( .B0(n5470), .B1(n4924), .A0N(n5125), .A1N(x_matrix[263]), 
        .Y(n4068) );
  OAI2BB2X1 U5960 ( .B0(n5492), .B1(n4924), .A0N(n5360), .A1N(x_matrix[359]), 
        .Y(n3940) );
  OAI2BB2X1 U5961 ( .B0(n5509), .B1(n4924), .A0N(n5141), .A1N(x_matrix[391]), 
        .Y(n3876) );
  OAI2BB2X1 U5962 ( .B0(n5514), .B1(n4924), .A0N(n5382), .A1N(x_matrix[455]), 
        .Y(n3812) );
  OAI2BB2X1 U5963 ( .B0(n5525), .B1(n4924), .A0N(n5151), .A1N(x_matrix[487]), 
        .Y(n3748) );
  OAI2BB2X1 U5964 ( .B0(n5407), .B1(n4923), .A0N(n5090), .A1N(x_matrix[8]), 
        .Y(n4451) );
  OAI2BB2X1 U5965 ( .B0(n5415), .B1(n4923), .A0N(n5343), .A1N(x_matrix[72]), 
        .Y(n4387) );
  OAI2BB2X1 U5966 ( .B0(n5429), .B1(n4923), .A0N(n5100), .A1N(x_matrix[88]), 
        .Y(n4323) );
  OAI2BB2X1 U5967 ( .B0(n5437), .B1(n4923), .A0N(n5356), .A1N(x_matrix[152]), 
        .Y(n4259) );
  OAI2BB2X1 U5968 ( .B0(n5448), .B1(n4923), .A0N(n5109), .A1N(x_matrix[168]), 
        .Y(n4195) );
  OAI2BB2X1 U5969 ( .B0(n5470), .B1(n4923), .A0N(n5125), .A1N(x_matrix[264]), 
        .Y(n4067) );
  OAI2BB2X1 U5970 ( .B0(n5492), .B1(n4923), .A0N(n5360), .A1N(x_matrix[360]), 
        .Y(n3939) );
  OAI2BB2X1 U5971 ( .B0(n5506), .B1(n4923), .A0N(n5142), .A1N(x_matrix[392]), 
        .Y(n3875) );
  OAI2BB2X1 U5972 ( .B0(n5514), .B1(n4923), .A0N(n5382), .A1N(x_matrix[456]), 
        .Y(n3811) );
  OAI2BB2X1 U5973 ( .B0(n5526), .B1(n4923), .A0N(n5151), .A1N(x_matrix[488]), 
        .Y(n3747) );
  OAI2BB2X1 U5974 ( .B0(n5409), .B1(n4922), .A0N(n5091), .A1N(x_matrix[9]), 
        .Y(n4450) );
  OAI2BB2X1 U5975 ( .B0(n5415), .B1(n4922), .A0N(n5341), .A1N(x_matrix[73]), 
        .Y(n4386) );
  OAI2BB2X1 U5976 ( .B0(n5431), .B1(n4922), .A0N(n5101), .A1N(x_matrix[89]), 
        .Y(n4322) );
  OAI2BB2X1 U5977 ( .B0(n5437), .B1(n4922), .A0N(n5354), .A1N(x_matrix[153]), 
        .Y(n4258) );
  OAI2BB2X1 U5978 ( .B0(n5448), .B1(n4922), .A0N(n5109), .A1N(x_matrix[169]), 
        .Y(n4194) );
  OAI2BB2X1 U5979 ( .B0(n5470), .B1(n4922), .A0N(n5125), .A1N(x_matrix[265]), 
        .Y(n4066) );
  OAI2BB2X1 U5980 ( .B0(n5492), .B1(n4922), .A0N(n5360), .A1N(x_matrix[361]), 
        .Y(n3938) );
  OAI2BB2X1 U5981 ( .B0(n5508), .B1(n4922), .A0N(n5143), .A1N(x_matrix[393]), 
        .Y(n3874) );
  OAI2BB2X1 U5982 ( .B0(n5514), .B1(n4922), .A0N(n5382), .A1N(x_matrix[457]), 
        .Y(n3810) );
  OAI2BB2X1 U5983 ( .B0(n5532), .B1(n4922), .A0N(n5151), .A1N(x_matrix[489]), 
        .Y(n3746) );
  OAI2BB2X1 U5984 ( .B0(n5404), .B1(n4978), .A0N(n5089), .A1N(x_matrix[16]), 
        .Y(n4443) );
  OAI2BB2X1 U5985 ( .B0(n5426), .B1(n4978), .A0N(n5099), .A1N(x_matrix[96]), 
        .Y(n4315) );
  OAI2BB2X1 U5986 ( .B0(n5449), .B1(n4978), .A0N(n5110), .A1N(x_matrix[176]), 
        .Y(n4187) );
  OAI2BB2X1 U5987 ( .B0(n5460), .B1(n4978), .A0N(n5117), .A1N(x_matrix[208]), 
        .Y(n4123) );
  OAI2BB2X1 U5988 ( .B0(n5471), .B1(n4978), .A0N(n5126), .A1N(x_matrix[272]), 
        .Y(n4059) );
  OAI2BB2X1 U5989 ( .B0(n5482), .B1(n4978), .A0N(n5133), .A1N(x_matrix[304]), 
        .Y(n3995) );
  OAI2BB2X1 U5990 ( .B0(n5503), .B1(n4978), .A0N(n5141), .A1N(x_matrix[400]), 
        .Y(n3867) );
  OAI2BB2X1 U5991 ( .B0(n5525), .B1(n4978), .A0N(n5152), .A1N(x_matrix[496]), 
        .Y(n3739) );
  OAI2BB2X1 U5992 ( .B0(n5537), .B1(n4978), .A0N(n5161), .A1N(x_matrix[544]), 
        .Y(n3675) );
  OAI2BB2X1 U5993 ( .B0(n5572), .B1(n4978), .A0N(n5169), .A1N(x_matrix[656]), 
        .Y(n3547) );
  OAI2BB2X1 U5994 ( .B0(n5404), .B1(n4977), .A0N(n5089), .A1N(x_matrix[17]), 
        .Y(n4442) );
  OAI2BB2X1 U5995 ( .B0(n5426), .B1(n4977), .A0N(n5099), .A1N(x_matrix[97]), 
        .Y(n4314) );
  OAI2BB2X1 U5996 ( .B0(n5449), .B1(n4977), .A0N(n5110), .A1N(x_matrix[177]), 
        .Y(n4186) );
  OAI2BB2X1 U5997 ( .B0(n5460), .B1(n4977), .A0N(n5117), .A1N(x_matrix[209]), 
        .Y(n4122) );
  OAI2BB2X1 U5998 ( .B0(n5471), .B1(n4977), .A0N(n5126), .A1N(x_matrix[273]), 
        .Y(n4058) );
  OAI2BB2X1 U5999 ( .B0(n5482), .B1(n4977), .A0N(n5134), .A1N(x_matrix[305]), 
        .Y(n3994) );
  OAI2BB2X1 U6000 ( .B0(n5503), .B1(n4977), .A0N(n5141), .A1N(x_matrix[401]), 
        .Y(n3866) );
  OAI2BB2X1 U6001 ( .B0(n5525), .B1(n4977), .A0N(n5152), .A1N(x_matrix[497]), 
        .Y(n3738) );
  OAI2BB2X1 U6002 ( .B0(n5537), .B1(n4977), .A0N(n5161), .A1N(x_matrix[545]), 
        .Y(n3674) );
  OAI2BB2X1 U6003 ( .B0(n5572), .B1(n4977), .A0N(n5169), .A1N(x_matrix[657]), 
        .Y(n3546) );
  OAI2BB2X1 U6004 ( .B0(n5404), .B1(n4976), .A0N(n5089), .A1N(x_matrix[18]), 
        .Y(n4441) );
  OAI2BB2X1 U6005 ( .B0(n5426), .B1(n4976), .A0N(n5099), .A1N(x_matrix[98]), 
        .Y(n4313) );
  OAI2BB2X1 U6006 ( .B0(n5449), .B1(n4976), .A0N(n5110), .A1N(x_matrix[178]), 
        .Y(n4185) );
  OAI2BB2X1 U6007 ( .B0(n5460), .B1(n4976), .A0N(n5117), .A1N(x_matrix[210]), 
        .Y(n4121) );
  OAI2BB2X1 U6008 ( .B0(n5471), .B1(n4976), .A0N(n5126), .A1N(x_matrix[274]), 
        .Y(n4057) );
  OAI2BB2X1 U6009 ( .B0(n5482), .B1(n4976), .A0N(n5135), .A1N(x_matrix[306]), 
        .Y(n3993) );
  OAI2BB2X1 U6010 ( .B0(n5503), .B1(n4976), .A0N(n5141), .A1N(x_matrix[402]), 
        .Y(n3865) );
  OAI2BB2X1 U6011 ( .B0(n5525), .B1(n4976), .A0N(n5152), .A1N(x_matrix[498]), 
        .Y(n3737) );
  OAI2BB2X1 U6012 ( .B0(n5537), .B1(n4976), .A0N(n5161), .A1N(x_matrix[546]), 
        .Y(n3673) );
  OAI2BB2X1 U6013 ( .B0(n5572), .B1(n4976), .A0N(n5169), .A1N(x_matrix[658]), 
        .Y(n3545) );
  OAI2BB2X1 U6014 ( .B0(n5404), .B1(n4975), .A0N(n5089), .A1N(x_matrix[19]), 
        .Y(n4440) );
  OAI2BB2X1 U6015 ( .B0(n5426), .B1(n4975), .A0N(n5099), .A1N(x_matrix[99]), 
        .Y(n4312) );
  OAI2BB2X1 U6016 ( .B0(n5449), .B1(n4975), .A0N(n5110), .A1N(x_matrix[179]), 
        .Y(n4184) );
  OAI2BB2X1 U6017 ( .B0(n5460), .B1(n4975), .A0N(n5117), .A1N(x_matrix[211]), 
        .Y(n4120) );
  OAI2BB2X1 U6018 ( .B0(n5471), .B1(n4975), .A0N(n5126), .A1N(x_matrix[275]), 
        .Y(n4056) );
  OAI2BB2X1 U6019 ( .B0(n5482), .B1(n4975), .A0N(n5133), .A1N(x_matrix[307]), 
        .Y(n3992) );
  OAI2BB2X1 U6020 ( .B0(n5503), .B1(n4975), .A0N(n5141), .A1N(x_matrix[403]), 
        .Y(n3864) );
  OAI2BB2X1 U6021 ( .B0(n5525), .B1(n4975), .A0N(n5152), .A1N(x_matrix[499]), 
        .Y(n3736) );
  OAI2BB2X1 U6022 ( .B0(n5537), .B1(n4975), .A0N(n5161), .A1N(x_matrix[547]), 
        .Y(n3672) );
  OAI2BB2X1 U6023 ( .B0(n5572), .B1(n4975), .A0N(n5169), .A1N(x_matrix[659]), 
        .Y(n3544) );
  OAI2BB2X1 U6024 ( .B0(n5404), .B1(n4973), .A0N(n5089), .A1N(x_matrix[20]), 
        .Y(n4439) );
  OAI2BB2X1 U6025 ( .B0(n5426), .B1(n4973), .A0N(n5099), .A1N(x_matrix[100]), 
        .Y(n4311) );
  OAI2BB2X1 U6026 ( .B0(n5449), .B1(n4973), .A0N(n5110), .A1N(x_matrix[180]), 
        .Y(n4183) );
  OAI2BB2X1 U6027 ( .B0(n5460), .B1(n4973), .A0N(n5117), .A1N(x_matrix[212]), 
        .Y(n4119) );
  OAI2BB2X1 U6028 ( .B0(n5471), .B1(n4973), .A0N(n5126), .A1N(x_matrix[276]), 
        .Y(n4055) );
  OAI2BB2X1 U6029 ( .B0(n5482), .B1(n4973), .A0N(n5134), .A1N(x_matrix[308]), 
        .Y(n3991) );
  OAI2BB2X1 U6030 ( .B0(n5503), .B1(n4973), .A0N(n5141), .A1N(x_matrix[404]), 
        .Y(n3863) );
  OAI2BB2X1 U6031 ( .B0(n5525), .B1(n4973), .A0N(n5152), .A1N(x_matrix[500]), 
        .Y(n3735) );
  OAI2BB2X1 U6032 ( .B0(n5537), .B1(n4973), .A0N(n5161), .A1N(x_matrix[548]), 
        .Y(n3671) );
  OAI2BB2X1 U6033 ( .B0(n5572), .B1(n4973), .A0N(n5169), .A1N(x_matrix[660]), 
        .Y(n3543) );
  OAI2BB2X1 U6034 ( .B0(n5404), .B1(n4972), .A0N(n5089), .A1N(x_matrix[21]), 
        .Y(n4438) );
  OAI2BB2X1 U6035 ( .B0(n5426), .B1(n4972), .A0N(n5099), .A1N(x_matrix[101]), 
        .Y(n4310) );
  OAI2BB2X1 U6036 ( .B0(n5449), .B1(n4972), .A0N(n5110), .A1N(x_matrix[181]), 
        .Y(n4182) );
  OAI2BB2X1 U6037 ( .B0(n5460), .B1(n4972), .A0N(n5117), .A1N(x_matrix[213]), 
        .Y(n4118) );
  OAI2BB2X1 U6038 ( .B0(n5471), .B1(n4972), .A0N(n5126), .A1N(x_matrix[277]), 
        .Y(n4054) );
  OAI2BB2X1 U6039 ( .B0(n5482), .B1(n4972), .A0N(n5135), .A1N(x_matrix[309]), 
        .Y(n3990) );
  OAI2BB2X1 U6040 ( .B0(n5503), .B1(n4972), .A0N(n5141), .A1N(x_matrix[405]), 
        .Y(n3862) );
  OAI2BB2X1 U6041 ( .B0(n5525), .B1(n4972), .A0N(n5152), .A1N(x_matrix[501]), 
        .Y(n3734) );
  OAI2BB2X1 U6042 ( .B0(n5537), .B1(n4972), .A0N(n5161), .A1N(x_matrix[549]), 
        .Y(n3670) );
  OAI2BB2X1 U6043 ( .B0(n5572), .B1(n4972), .A0N(n5169), .A1N(x_matrix[661]), 
        .Y(n3542) );
  OAI2BB2X1 U6044 ( .B0(n5404), .B1(n4971), .A0N(n5089), .A1N(x_matrix[22]), 
        .Y(n4437) );
  OAI2BB2X1 U6045 ( .B0(n5426), .B1(n4971), .A0N(n5099), .A1N(x_matrix[102]), 
        .Y(n4309) );
  OAI2BB2X1 U6046 ( .B0(n5449), .B1(n4971), .A0N(n5110), .A1N(x_matrix[182]), 
        .Y(n4181) );
  OAI2BB2X1 U6047 ( .B0(n5460), .B1(n4971), .A0N(n5117), .A1N(x_matrix[214]), 
        .Y(n4117) );
  OAI2BB2X1 U6048 ( .B0(n5471), .B1(n4971), .A0N(n5126), .A1N(x_matrix[278]), 
        .Y(n4053) );
  OAI2BB2X1 U6049 ( .B0(n5482), .B1(n4971), .A0N(n5133), .A1N(x_matrix[310]), 
        .Y(n3989) );
  OAI2BB2X1 U6050 ( .B0(n5503), .B1(n4971), .A0N(n5141), .A1N(x_matrix[406]), 
        .Y(n3861) );
  OAI2BB2X1 U6051 ( .B0(n5525), .B1(n4971), .A0N(n5152), .A1N(x_matrix[502]), 
        .Y(n3733) );
  OAI2BB2X1 U6052 ( .B0(n5537), .B1(n4971), .A0N(n5161), .A1N(x_matrix[550]), 
        .Y(n3669) );
  OAI2BB2X1 U6053 ( .B0(n5572), .B1(n4971), .A0N(n5169), .A1N(x_matrix[662]), 
        .Y(n3541) );
  OAI2BB2X1 U6054 ( .B0(n5404), .B1(n4970), .A0N(n5089), .A1N(x_matrix[23]), 
        .Y(n4436) );
  OAI2BB2X1 U6055 ( .B0(n5426), .B1(n4970), .A0N(n5099), .A1N(x_matrix[103]), 
        .Y(n4308) );
  OAI2BB2X1 U6056 ( .B0(n5449), .B1(n4970), .A0N(n5110), .A1N(x_matrix[183]), 
        .Y(n4180) );
  OAI2BB2X1 U6057 ( .B0(n5460), .B1(n4970), .A0N(n5117), .A1N(x_matrix[215]), 
        .Y(n4116) );
  OAI2BB2X1 U6058 ( .B0(n5471), .B1(n4970), .A0N(n5126), .A1N(x_matrix[279]), 
        .Y(n4052) );
  OAI2BB2X1 U6059 ( .B0(n5482), .B1(n4970), .A0N(n5134), .A1N(x_matrix[311]), 
        .Y(n3988) );
  OAI2BB2X1 U6060 ( .B0(n5503), .B1(n4970), .A0N(n5141), .A1N(x_matrix[407]), 
        .Y(n3860) );
  OAI2BB2X1 U6061 ( .B0(n5525), .B1(n4970), .A0N(n5152), .A1N(x_matrix[503]), 
        .Y(n3732) );
  OAI2BB2X1 U6062 ( .B0(n5537), .B1(n4970), .A0N(n5161), .A1N(x_matrix[551]), 
        .Y(n3668) );
  OAI2BB2X1 U6063 ( .B0(n5572), .B1(n4970), .A0N(n5169), .A1N(x_matrix[663]), 
        .Y(n3540) );
  OAI2BB2X1 U6064 ( .B0(n5404), .B1(n4969), .A0N(n5090), .A1N(x_matrix[24]), 
        .Y(n4435) );
  OAI2BB2X1 U6065 ( .B0(n5426), .B1(n4969), .A0N(n5100), .A1N(x_matrix[104]), 
        .Y(n4307) );
  OAI2BB2X1 U6066 ( .B0(n5449), .B1(n4969), .A0N(n5111), .A1N(x_matrix[184]), 
        .Y(n4179) );
  OAI2BB2X1 U6067 ( .B0(n5460), .B1(n4969), .A0N(n5117), .A1N(x_matrix[216]), 
        .Y(n4115) );
  OAI2BB2X1 U6068 ( .B0(n5471), .B1(n4969), .A0N(n5127), .A1N(x_matrix[280]), 
        .Y(n4051) );
  OAI2BB2X1 U6069 ( .B0(n5482), .B1(n4969), .A0N(n5135), .A1N(x_matrix[312]), 
        .Y(n3987) );
  OAI2BB2X1 U6070 ( .B0(n5503), .B1(n4969), .A0N(n5142), .A1N(x_matrix[408]), 
        .Y(n3859) );
  OAI2BB2X1 U6071 ( .B0(n5526), .B1(n4969), .A0N(n5153), .A1N(x_matrix[504]), 
        .Y(n3731) );
  OAI2BB2X1 U6072 ( .B0(n5537), .B1(n4969), .A0N(n5161), .A1N(x_matrix[552]), 
        .Y(n3667) );
  OAI2BB2X1 U6073 ( .B0(n5572), .B1(n4969), .A0N(n5169), .A1N(x_matrix[664]), 
        .Y(n3539) );
  OAI2BB2X1 U6074 ( .B0(n5404), .B1(n4968), .A0N(n5090), .A1N(x_matrix[25]), 
        .Y(n4434) );
  OAI2BB2X1 U6075 ( .B0(n5426), .B1(n4968), .A0N(n5100), .A1N(x_matrix[105]), 
        .Y(n4306) );
  OAI2BB2X1 U6076 ( .B0(n5454), .B1(n4968), .A0N(n5111), .A1N(x_matrix[185]), 
        .Y(n4178) );
  OAI2BB2X1 U6077 ( .B0(n5460), .B1(n4968), .A0N(n5117), .A1N(x_matrix[217]), 
        .Y(n4114) );
  OAI2BB2X1 U6078 ( .B0(n5476), .B1(n4968), .A0N(n5127), .A1N(x_matrix[281]), 
        .Y(n4050) );
  OAI2BB2X1 U6079 ( .B0(n5482), .B1(n4968), .A0N(n5140), .A1N(x_matrix[313]), 
        .Y(n3986) );
  OAI2BB2X1 U6080 ( .B0(n5503), .B1(n4968), .A0N(n5142), .A1N(x_matrix[409]), 
        .Y(n3858) );
  OAI2BB2X1 U6081 ( .B0(n5526), .B1(n4968), .A0N(n5153), .A1N(x_matrix[505]), 
        .Y(n3730) );
  OAI2BB2X1 U6082 ( .B0(n5537), .B1(n4968), .A0N(n5161), .A1N(x_matrix[553]), 
        .Y(n3666) );
  OAI2BB2X1 U6083 ( .B0(n5572), .B1(n4968), .A0N(n5169), .A1N(x_matrix[665]), 
        .Y(n3538) );
  OAI2BB2X1 U6084 ( .B0(n5404), .B1(n4967), .A0N(n5090), .A1N(x_matrix[26]), 
        .Y(n4433) );
  OAI2BB2X1 U6085 ( .B0(n5426), .B1(n4967), .A0N(n5100), .A1N(x_matrix[106]), 
        .Y(n4305) );
  OAI2BB2X1 U6086 ( .B0(n5449), .B1(n4967), .A0N(n5111), .A1N(x_matrix[186]), 
        .Y(n4177) );
  OAI2BB2X1 U6087 ( .B0(n5460), .B1(n4967), .A0N(n5117), .A1N(x_matrix[218]), 
        .Y(n4113) );
  OAI2BB2X1 U6088 ( .B0(n5471), .B1(n4967), .A0N(n5127), .A1N(x_matrix[282]), 
        .Y(n4049) );
  OAI2BB2X1 U6089 ( .B0(n5482), .B1(n4967), .A0N(n5133), .A1N(x_matrix[314]), 
        .Y(n3985) );
  OAI2BB2X1 U6090 ( .B0(n5503), .B1(n4967), .A0N(n5142), .A1N(x_matrix[410]), 
        .Y(n3857) );
  OAI2BB2X1 U6091 ( .B0(n5526), .B1(n4967), .A0N(n5153), .A1N(x_matrix[506]), 
        .Y(n3729) );
  OAI2BB2X1 U6092 ( .B0(n5537), .B1(n4967), .A0N(n5161), .A1N(x_matrix[554]), 
        .Y(n3665) );
  OAI2BB2X1 U6093 ( .B0(n5572), .B1(n4967), .A0N(n5169), .A1N(x_matrix[666]), 
        .Y(n3537) );
  OAI2BB2X1 U6094 ( .B0(n5404), .B1(n4966), .A0N(n5090), .A1N(x_matrix[27]), 
        .Y(n4432) );
  OAI2BB2X1 U6095 ( .B0(n5426), .B1(n4966), .A0N(n5100), .A1N(x_matrix[107]), 
        .Y(n4304) );
  OAI2BB2X1 U6096 ( .B0(n5454), .B1(n4966), .A0N(n5111), .A1N(x_matrix[187]), 
        .Y(n4176) );
  OAI2BB2X1 U6097 ( .B0(n5460), .B1(n4966), .A0N(n5117), .A1N(x_matrix[219]), 
        .Y(n4112) );
  OAI2BB2X1 U6098 ( .B0(n5476), .B1(n4966), .A0N(n5127), .A1N(x_matrix[283]), 
        .Y(n4048) );
  OAI2BB2X1 U6099 ( .B0(n5482), .B1(n4966), .A0N(n5134), .A1N(x_matrix[315]), 
        .Y(n3984) );
  OAI2BB2X1 U6100 ( .B0(n5503), .B1(n4966), .A0N(n5142), .A1N(x_matrix[411]), 
        .Y(n3856) );
  OAI2BB2X1 U6101 ( .B0(n5526), .B1(n4966), .A0N(n5153), .A1N(x_matrix[507]), 
        .Y(n3728) );
  OAI2BB2X1 U6102 ( .B0(n5537), .B1(n4966), .A0N(n5161), .A1N(x_matrix[555]), 
        .Y(n3664) );
  OAI2BB2X1 U6103 ( .B0(n5572), .B1(n4966), .A0N(n5169), .A1N(x_matrix[667]), 
        .Y(n3536) );
  OAI2BB2X1 U6104 ( .B0(n5405), .B1(n4965), .A0N(n5090), .A1N(x_matrix[28]), 
        .Y(n4431) );
  OAI2BB2X1 U6105 ( .B0(n5427), .B1(n4965), .A0N(n5100), .A1N(x_matrix[108]), 
        .Y(n4303) );
  OAI2BB2X1 U6106 ( .B0(n5449), .B1(n4965), .A0N(n5111), .A1N(x_matrix[188]), 
        .Y(n4175) );
  OAI2BB2X1 U6107 ( .B0(n5459), .B1(n4965), .A0N(n5118), .A1N(x_matrix[220]), 
        .Y(n4111) );
  OAI2BB2X1 U6108 ( .B0(n5471), .B1(n4965), .A0N(n5127), .A1N(x_matrix[284]), 
        .Y(n4047) );
  OAI2BB2X1 U6109 ( .B0(n5481), .B1(n4965), .A0N(n5133), .A1N(x_matrix[316]), 
        .Y(n3983) );
  OAI2BB2X1 U6110 ( .B0(n5504), .B1(n4965), .A0N(n5142), .A1N(x_matrix[412]), 
        .Y(n3855) );
  OAI2BB2X1 U6111 ( .B0(n5526), .B1(n4965), .A0N(n5153), .A1N(x_matrix[508]), 
        .Y(n3727) );
  OAI2BB2X1 U6112 ( .B0(n5536), .B1(n4965), .A0N(n5162), .A1N(x_matrix[556]), 
        .Y(n3663) );
  OAI2BB2X1 U6113 ( .B0(n5571), .B1(n4965), .A0N(n5170), .A1N(x_matrix[668]), 
        .Y(n3535) );
  OAI2BB2X1 U6114 ( .B0(n5406), .B1(n4964), .A0N(n5090), .A1N(x_matrix[29]), 
        .Y(n4430) );
  OAI2BB2X1 U6115 ( .B0(n5428), .B1(n4964), .A0N(n5100), .A1N(x_matrix[109]), 
        .Y(n4302) );
  OAI2BB2X1 U6116 ( .B0(n5454), .B1(n4964), .A0N(n5111), .A1N(x_matrix[189]), 
        .Y(n4174) );
  OAI2BB2X1 U6117 ( .B0(n5459), .B1(n4964), .A0N(n5118), .A1N(x_matrix[221]), 
        .Y(n4110) );
  OAI2BB2X1 U6118 ( .B0(n5476), .B1(n4964), .A0N(n5127), .A1N(x_matrix[285]), 
        .Y(n4046) );
  OAI2BB2X1 U6119 ( .B0(n5481), .B1(n4964), .A0N(n5133), .A1N(x_matrix[317]), 
        .Y(n3982) );
  OAI2BB2X1 U6120 ( .B0(n5505), .B1(n4964), .A0N(n5142), .A1N(x_matrix[413]), 
        .Y(n3854) );
  OAI2BB2X1 U6121 ( .B0(n5526), .B1(n4964), .A0N(n5153), .A1N(x_matrix[509]), 
        .Y(n3726) );
  OAI2BB2X1 U6122 ( .B0(n5536), .B1(n4964), .A0N(n5162), .A1N(x_matrix[557]), 
        .Y(n3662) );
  OAI2BB2X1 U6123 ( .B0(n5571), .B1(n4964), .A0N(n5170), .A1N(x_matrix[669]), 
        .Y(n3534) );
  OAI2BB2X1 U6124 ( .B0(n5405), .B1(n4962), .A0N(n5090), .A1N(x_matrix[30]), 
        .Y(n4429) );
  OAI2BB2X1 U6125 ( .B0(n5427), .B1(n4962), .A0N(n5100), .A1N(x_matrix[110]), 
        .Y(n4301) );
  OAI2BB2X1 U6126 ( .B0(n5449), .B1(n4962), .A0N(n5111), .A1N(x_matrix[190]), 
        .Y(n4173) );
  OAI2BB2X1 U6127 ( .B0(n5459), .B1(n4962), .A0N(n5118), .A1N(x_matrix[222]), 
        .Y(n4109) );
  OAI2BB2X1 U6128 ( .B0(n5471), .B1(n4962), .A0N(n5127), .A1N(x_matrix[286]), 
        .Y(n4045) );
  OAI2BB2X1 U6129 ( .B0(n5481), .B1(n4962), .A0N(n5133), .A1N(x_matrix[318]), 
        .Y(n3981) );
  OAI2BB2X1 U6130 ( .B0(n5504), .B1(n4962), .A0N(n5142), .A1N(x_matrix[414]), 
        .Y(n3853) );
  OAI2BB2X1 U6131 ( .B0(n5526), .B1(n4962), .A0N(n5153), .A1N(x_matrix[510]), 
        .Y(n3725) );
  OAI2BB2X1 U6132 ( .B0(n5536), .B1(n4962), .A0N(n5162), .A1N(x_matrix[558]), 
        .Y(n3661) );
  OAI2BB2X1 U6133 ( .B0(n5571), .B1(n4962), .A0N(n5170), .A1N(x_matrix[670]), 
        .Y(n3533) );
  OAI2BB2X1 U6134 ( .B0(n5406), .B1(n4961), .A0N(n5090), .A1N(x_matrix[31]), 
        .Y(n4428) );
  OAI2BB2X1 U6135 ( .B0(n5428), .B1(n4961), .A0N(n5100), .A1N(x_matrix[111]), 
        .Y(n4300) );
  OAI2BB2X1 U6136 ( .B0(n5454), .B1(n4961), .A0N(n5111), .A1N(x_matrix[191]), 
        .Y(n4172) );
  OAI2BB2X1 U6137 ( .B0(n5459), .B1(n4961), .A0N(n5118), .A1N(x_matrix[223]), 
        .Y(n4108) );
  OAI2BB2X1 U6138 ( .B0(n5476), .B1(n4961), .A0N(n5127), .A1N(x_matrix[287]), 
        .Y(n4044) );
  OAI2BB2X1 U6139 ( .B0(n5481), .B1(n4961), .A0N(n5133), .A1N(x_matrix[319]), 
        .Y(n3980) );
  OAI2BB2X1 U6140 ( .B0(n5505), .B1(n4961), .A0N(n5142), .A1N(x_matrix[415]), 
        .Y(n3852) );
  OAI2BB2X1 U6141 ( .B0(n5526), .B1(n4961), .A0N(n5153), .A1N(x_matrix[511]), 
        .Y(n3724) );
  OAI2BB2X1 U6142 ( .B0(n5536), .B1(n4961), .A0N(n5162), .A1N(x_matrix[559]), 
        .Y(n3660) );
  OAI2BB2X1 U6143 ( .B0(n5571), .B1(n4961), .A0N(n5170), .A1N(x_matrix[671]), 
        .Y(n3532) );
  OAI2BB2X1 U6144 ( .B0(n5406), .B1(n4943), .A0N(n5092), .A1N(x_matrix[48]), 
        .Y(n4411) );
  OAI2BB2X1 U6145 ( .B0(n5428), .B1(n4943), .A0N(n5102), .A1N(x_matrix[128]), 
        .Y(n4283) );
  OAI2BB2X1 U6146 ( .B0(n5459), .B1(n4943), .A0N(n5119), .A1N(x_matrix[240]), 
        .Y(n4091) );
  OAI2BB2X1 U6147 ( .B0(n5481), .B1(n4943), .A0N(n5134), .A1N(x_matrix[336]), 
        .Y(n3963) );
  OAI2BB2X1 U6148 ( .B0(n5494), .B1(n4943), .A0N(n5361), .A1N(x_matrix[368]), 
        .Y(n3899) );
  OAI2BB2X1 U6149 ( .B0(n5505), .B1(n4943), .A0N(n5144), .A1N(x_matrix[432]), 
        .Y(n3835) );
  OAI2BB2X1 U6150 ( .B0(n5516), .B1(n4943), .A0N(n5383), .A1N(x_matrix[464]), 
        .Y(n3771) );
  OAI2BB2X1 U6151 ( .B0(n5528), .B1(n4943), .A0N(n5154), .A1N(x_matrix[528]), 
        .Y(n3707) );
  OAI2BB2X1 U6152 ( .B0(n5536), .B1(n4943), .A0N(n5163), .A1N(x_matrix[576]), 
        .Y(n3643) );
  OAI2BB2X1 U6153 ( .B0(n5571), .B1(n4943), .A0N(n5171), .A1N(x_matrix[688]), 
        .Y(n3515) );
  OAI2BB2X1 U6154 ( .B0(n5406), .B1(n4942), .A0N(n5097), .A1N(x_matrix[49]), 
        .Y(n4410) );
  OAI2BB2X1 U6155 ( .B0(n5428), .B1(n4942), .A0N(n5107), .A1N(x_matrix[129]), 
        .Y(n4282) );
  OAI2BB2X1 U6156 ( .B0(n5465), .B1(n4942), .A0N(n5119), .A1N(x_matrix[241]), 
        .Y(n4090) );
  OAI2BB2X1 U6157 ( .B0(n5487), .B1(n4942), .A0N(n5134), .A1N(x_matrix[337]), 
        .Y(n3962) );
  OAI2BB2X1 U6158 ( .B0(n5493), .B1(n4942), .A0N(n5361), .A1N(x_matrix[369]), 
        .Y(n3898) );
  OAI2BB2X1 U6159 ( .B0(n5505), .B1(n4942), .A0N(n5149), .A1N(x_matrix[433]), 
        .Y(n3834) );
  OAI2BB2X1 U6160 ( .B0(n5515), .B1(n4942), .A0N(n5383), .A1N(x_matrix[465]), 
        .Y(n3770) );
  OAI2BB2X1 U6161 ( .B0(n5528), .B1(n4942), .A0N(n5154), .A1N(x_matrix[529]), 
        .Y(n3706) );
  OAI2BB2X1 U6162 ( .B0(n5542), .B1(n4942), .A0N(n5163), .A1N(x_matrix[577]), 
        .Y(n3642) );
  OAI2BB2X1 U6163 ( .B0(n5577), .B1(n4942), .A0N(n5171), .A1N(x_matrix[689]), 
        .Y(n3514) );
  OAI2BB2X1 U6164 ( .B0(n5406), .B1(n4940), .A0N(n5091), .A1N(x_matrix[50]), 
        .Y(n4409) );
  OAI2BB2X1 U6165 ( .B0(n5428), .B1(n4940), .A0N(n5101), .A1N(x_matrix[130]), 
        .Y(n4281) );
  OAI2BB2X1 U6166 ( .B0(n5459), .B1(n4940), .A0N(n5119), .A1N(x_matrix[242]), 
        .Y(n4089) );
  OAI2BB2X1 U6167 ( .B0(n5481), .B1(n4940), .A0N(n5134), .A1N(x_matrix[338]), 
        .Y(n3961) );
  OAI2BB2X1 U6168 ( .B0(n5493), .B1(n4940), .A0N(n5361), .A1N(x_matrix[370]), 
        .Y(n3897) );
  OAI2BB2X1 U6169 ( .B0(n5505), .B1(n4940), .A0N(n5143), .A1N(x_matrix[434]), 
        .Y(n3833) );
  OAI2BB2X1 U6170 ( .B0(n5515), .B1(n4940), .A0N(n5383), .A1N(x_matrix[466]), 
        .Y(n3769) );
  OAI2BB2X1 U6171 ( .B0(n5528), .B1(n4940), .A0N(n5154), .A1N(x_matrix[530]), 
        .Y(n3705) );
  OAI2BB2X1 U6172 ( .B0(n5536), .B1(n4940), .A0N(n5163), .A1N(x_matrix[578]), 
        .Y(n3641) );
  OAI2BB2X1 U6173 ( .B0(n5571), .B1(n4940), .A0N(n5171), .A1N(x_matrix[690]), 
        .Y(n3513) );
  OAI2BB2X1 U6174 ( .B0(n5406), .B1(n4939), .A0N(n5090), .A1N(x_matrix[51]), 
        .Y(n4408) );
  OAI2BB2X1 U6175 ( .B0(n5428), .B1(n4939), .A0N(n5100), .A1N(x_matrix[131]), 
        .Y(n4280) );
  OAI2BB2X1 U6176 ( .B0(n5465), .B1(n4939), .A0N(n5119), .A1N(x_matrix[243]), 
        .Y(n4088) );
  OAI2BB2X1 U6177 ( .B0(n5487), .B1(n4939), .A0N(n5134), .A1N(x_matrix[339]), 
        .Y(n3960) );
  OAI2BB2X1 U6178 ( .B0(n5493), .B1(n4939), .A0N(n5361), .A1N(x_matrix[371]), 
        .Y(n3896) );
  OAI2BB2X1 U6179 ( .B0(n5505), .B1(n4939), .A0N(n5142), .A1N(x_matrix[435]), 
        .Y(n3832) );
  OAI2BB2X1 U6180 ( .B0(n5515), .B1(n4939), .A0N(n5383), .A1N(x_matrix[467]), 
        .Y(n3768) );
  OAI2BB2X1 U6181 ( .B0(n5528), .B1(n4939), .A0N(n5154), .A1N(x_matrix[531]), 
        .Y(n3704) );
  OAI2BB2X1 U6182 ( .B0(n5542), .B1(n4939), .A0N(n5163), .A1N(x_matrix[579]), 
        .Y(n3640) );
  OAI2BB2X1 U6183 ( .B0(n5577), .B1(n4939), .A0N(n5171), .A1N(x_matrix[691]), 
        .Y(n3512) );
  OAI2BB2X1 U6184 ( .B0(n5406), .B1(n4938), .A0N(n5089), .A1N(x_matrix[52]), 
        .Y(n4407) );
  OAI2BB2X1 U6185 ( .B0(n5428), .B1(n4938), .A0N(n5099), .A1N(x_matrix[132]), 
        .Y(n4279) );
  OAI2BB2X1 U6186 ( .B0(n5466), .B1(n4938), .A0N(n5119), .A1N(x_matrix[244]), 
        .Y(n4087) );
  OAI2BB2X1 U6187 ( .B0(n5488), .B1(n4938), .A0N(n5135), .A1N(x_matrix[340]), 
        .Y(n3959) );
  OAI2BB2X1 U6188 ( .B0(n5497), .B1(n4938), .A0N(n5361), .A1N(x_matrix[372]), 
        .Y(n3895) );
  OAI2BB2X1 U6189 ( .B0(n5505), .B1(n4938), .A0N(n5141), .A1N(x_matrix[436]), 
        .Y(n3831) );
  OAI2BB2X1 U6190 ( .B0(n5519), .B1(n4938), .A0N(n5383), .A1N(x_matrix[468]), 
        .Y(n3767) );
  OAI2BB2X1 U6191 ( .B0(n5528), .B1(n4938), .A0N(n5154), .A1N(x_matrix[532]), 
        .Y(n3703) );
  OAI2BB2X1 U6192 ( .B0(n5543), .B1(n4938), .A0N(n5163), .A1N(x_matrix[580]), 
        .Y(n3639) );
  OAI2BB2X1 U6193 ( .B0(n5578), .B1(n4938), .A0N(n5171), .A1N(x_matrix[692]), 
        .Y(n3511) );
  OAI2BB2X1 U6194 ( .B0(n5406), .B1(n4937), .A0N(n5097), .A1N(x_matrix[53]), 
        .Y(n4406) );
  OAI2BB2X1 U6195 ( .B0(n5428), .B1(n4937), .A0N(n5107), .A1N(x_matrix[133]), 
        .Y(n4278) );
  OAI2BB2X1 U6196 ( .B0(n5466), .B1(n4937), .A0N(n5119), .A1N(x_matrix[245]), 
        .Y(n4086) );
  OAI2BB2X1 U6197 ( .B0(n5488), .B1(n4937), .A0N(n5135), .A1N(x_matrix[341]), 
        .Y(n3958) );
  OAI2BB2X1 U6198 ( .B0(n5493), .B1(n4937), .A0N(n5361), .A1N(x_matrix[373]), 
        .Y(n3894) );
  OAI2BB2X1 U6199 ( .B0(n5505), .B1(n4937), .A0N(n5149), .A1N(x_matrix[437]), 
        .Y(n3830) );
  OAI2BB2X1 U6200 ( .B0(n5515), .B1(n4937), .A0N(n5383), .A1N(x_matrix[469]), 
        .Y(n3766) );
  OAI2BB2X1 U6201 ( .B0(n5528), .B1(n4937), .A0N(n5154), .A1N(x_matrix[533]), 
        .Y(n3702) );
  OAI2BB2X1 U6202 ( .B0(n5543), .B1(n4937), .A0N(n5163), .A1N(x_matrix[581]), 
        .Y(n3638) );
  OAI2BB2X1 U6203 ( .B0(n5578), .B1(n4937), .A0N(n5171), .A1N(x_matrix[693]), 
        .Y(n3510) );
  OAI2BB2X1 U6204 ( .B0(n5406), .B1(n4936), .A0N(n5091), .A1N(x_matrix[54]), 
        .Y(n4405) );
  OAI2BB2X1 U6205 ( .B0(n5428), .B1(n4936), .A0N(n5101), .A1N(x_matrix[134]), 
        .Y(n4277) );
  OAI2BB2X1 U6206 ( .B0(n5460), .B1(n4936), .A0N(n5119), .A1N(x_matrix[246]), 
        .Y(n4085) );
  OAI2BB2X1 U6207 ( .B0(n5482), .B1(n4936), .A0N(n5135), .A1N(x_matrix[342]), 
        .Y(n3957) );
  OAI2BB2X1 U6208 ( .B0(n5499), .B1(n4936), .A0N(n5361), .A1N(x_matrix[374]), 
        .Y(n3893) );
  OAI2BB2X1 U6209 ( .B0(n5505), .B1(n4936), .A0N(n5143), .A1N(x_matrix[438]), 
        .Y(n3829) );
  OAI2BB2X1 U6210 ( .B0(n5521), .B1(n4936), .A0N(n5383), .A1N(x_matrix[470]), 
        .Y(n3765) );
  OAI2BB2X1 U6211 ( .B0(n5528), .B1(n4936), .A0N(n5154), .A1N(x_matrix[534]), 
        .Y(n3701) );
  OAI2BB2X1 U6212 ( .B0(n5537), .B1(n4936), .A0N(n5163), .A1N(x_matrix[582]), 
        .Y(n3637) );
  OAI2BB2X1 U6213 ( .B0(n5572), .B1(n4936), .A0N(n5171), .A1N(x_matrix[694]), 
        .Y(n3509) );
  OAI2BB2X1 U6214 ( .B0(n5406), .B1(n4935), .A0N(n5090), .A1N(x_matrix[55]), 
        .Y(n4404) );
  OAI2BB2X1 U6215 ( .B0(n5428), .B1(n4935), .A0N(n5100), .A1N(x_matrix[135]), 
        .Y(n4276) );
  OAI2BB2X1 U6216 ( .B0(n5460), .B1(n4935), .A0N(n5119), .A1N(x_matrix[247]), 
        .Y(n4084) );
  OAI2BB2X1 U6217 ( .B0(n5482), .B1(n4935), .A0N(n5135), .A1N(x_matrix[343]), 
        .Y(n3956) );
  OAI2BB2X1 U6218 ( .B0(n5493), .B1(n4935), .A0N(n5361), .A1N(x_matrix[375]), 
        .Y(n3892) );
  OAI2BB2X1 U6219 ( .B0(n5505), .B1(n4935), .A0N(n5142), .A1N(x_matrix[439]), 
        .Y(n3828) );
  OAI2BB2X1 U6220 ( .B0(n5515), .B1(n4935), .A0N(n5383), .A1N(x_matrix[471]), 
        .Y(n3764) );
  OAI2BB2X1 U6221 ( .B0(n5528), .B1(n4935), .A0N(n5154), .A1N(x_matrix[535]), 
        .Y(n3700) );
  OAI2BB2X1 U6222 ( .B0(n5537), .B1(n4935), .A0N(n5163), .A1N(x_matrix[583]), 
        .Y(n3636) );
  OAI2BB2X1 U6223 ( .B0(n5572), .B1(n4935), .A0N(n5171), .A1N(x_matrix[695]), 
        .Y(n3508) );
  OAI2BB2X1 U6224 ( .B0(n5406), .B1(n4934), .A0N(n5089), .A1N(x_matrix[56]), 
        .Y(n4403) );
  OAI2BB2X1 U6225 ( .B0(n5428), .B1(n4934), .A0N(n5099), .A1N(x_matrix[136]), 
        .Y(n4275) );
  OAI2BB2X1 U6226 ( .B0(n5461), .B1(n4934), .A0N(n5119), .A1N(x_matrix[248]), 
        .Y(n4083) );
  OAI2BB2X1 U6227 ( .B0(n5483), .B1(n4934), .A0N(n5135), .A1N(x_matrix[344]), 
        .Y(n3955) );
  OAI2BB2X1 U6228 ( .B0(n5498), .B1(n4934), .A0N(n5362), .A1N(x_matrix[376]), 
        .Y(n3891) );
  OAI2BB2X1 U6229 ( .B0(n5505), .B1(n4934), .A0N(n5141), .A1N(x_matrix[440]), 
        .Y(n3827) );
  OAI2BB2X1 U6230 ( .B0(n5520), .B1(n4934), .A0N(n5384), .A1N(x_matrix[472]), 
        .Y(n3763) );
  OAI2BB2X1 U6231 ( .B0(n5528), .B1(n4934), .A0N(n5154), .A1N(x_matrix[536]), 
        .Y(n3699) );
  OAI2BB2X1 U6232 ( .B0(n5538), .B1(n4934), .A0N(n5163), .A1N(x_matrix[584]), 
        .Y(n3635) );
  OAI2BB2X1 U6233 ( .B0(n5573), .B1(n4934), .A0N(n5171), .A1N(x_matrix[696]), 
        .Y(n3507) );
  OAI2BB2X1 U6234 ( .B0(n5406), .B1(n4933), .A0N(n5097), .A1N(x_matrix[57]), 
        .Y(n4402) );
  OAI2BB2X1 U6235 ( .B0(n5428), .B1(n4933), .A0N(n5107), .A1N(x_matrix[137]), 
        .Y(n4274) );
  OAI2BB2X1 U6236 ( .B0(n5460), .B1(n4933), .A0N(n5119), .A1N(x_matrix[249]), 
        .Y(n4082) );
  OAI2BB2X1 U6237 ( .B0(n5482), .B1(n4933), .A0N(n5135), .A1N(x_matrix[345]), 
        .Y(n3954) );
  OAI2BB2X1 U6238 ( .B0(n5493), .B1(n4933), .A0N(n5362), .A1N(x_matrix[377]), 
        .Y(n3890) );
  OAI2BB2X1 U6239 ( .B0(n5505), .B1(n4933), .A0N(n5149), .A1N(x_matrix[441]), 
        .Y(n3826) );
  OAI2BB2X1 U6240 ( .B0(n5515), .B1(n4933), .A0N(n5384), .A1N(x_matrix[473]), 
        .Y(n3762) );
  OAI2BB2X1 U6241 ( .B0(n5528), .B1(n4933), .A0N(n5154), .A1N(x_matrix[537]), 
        .Y(n3698) );
  OAI2BB2X1 U6242 ( .B0(n5537), .B1(n4933), .A0N(n5163), .A1N(x_matrix[585]), 
        .Y(n3634) );
  OAI2BB2X1 U6243 ( .B0(n5572), .B1(n4933), .A0N(n5171), .A1N(x_matrix[697]), 
        .Y(n3506) );
  OAI2BB2X1 U6244 ( .B0(n5406), .B1(n4932), .A0N(n5091), .A1N(x_matrix[58]), 
        .Y(n4401) );
  OAI2BB2X1 U6245 ( .B0(n5428), .B1(n4932), .A0N(n5101), .A1N(x_matrix[138]), 
        .Y(n4273) );
  OAI2BB2X1 U6246 ( .B0(n5461), .B1(n4932), .A0N(n5119), .A1N(x_matrix[250]), 
        .Y(n4081) );
  OAI2BB2X1 U6247 ( .B0(n5483), .B1(n4932), .A0N(n5135), .A1N(x_matrix[346]), 
        .Y(n3953) );
  OAI2BB2X1 U6248 ( .B0(n5492), .B1(n4932), .A0N(n5362), .A1N(x_matrix[378]), 
        .Y(n3889) );
  OAI2BB2X1 U6249 ( .B0(n5505), .B1(n4932), .A0N(n5143), .A1N(x_matrix[442]), 
        .Y(n3825) );
  OAI2BB2X1 U6250 ( .B0(n5514), .B1(n4932), .A0N(n5384), .A1N(x_matrix[474]), 
        .Y(n3761) );
  OAI2BB2X1 U6251 ( .B0(n5528), .B1(n4932), .A0N(n5154), .A1N(x_matrix[538]), 
        .Y(n3697) );
  OAI2BB2X1 U6252 ( .B0(n5538), .B1(n4932), .A0N(n5163), .A1N(x_matrix[586]), 
        .Y(n3633) );
  OAI2BB2X1 U6253 ( .B0(n5573), .B1(n4932), .A0N(n5171), .A1N(x_matrix[698]), 
        .Y(n3505) );
  OAI2BB2X1 U6254 ( .B0(n5406), .B1(n4931), .A0N(n5090), .A1N(x_matrix[59]), 
        .Y(n4400) );
  OAI2BB2X1 U6255 ( .B0(n5428), .B1(n4931), .A0N(n5100), .A1N(x_matrix[139]), 
        .Y(n4272) );
  OAI2BB2X1 U6256 ( .B0(n5460), .B1(n4931), .A0N(n5119), .A1N(x_matrix[251]), 
        .Y(n4080) );
  OAI2BB2X1 U6257 ( .B0(n5482), .B1(n4931), .A0N(n5135), .A1N(x_matrix[347]), 
        .Y(n3952) );
  OAI2BB2X1 U6258 ( .B0(n5493), .B1(n4931), .A0N(n5362), .A1N(x_matrix[379]), 
        .Y(n3888) );
  OAI2BB2X1 U6259 ( .B0(n5505), .B1(n4931), .A0N(n5142), .A1N(x_matrix[443]), 
        .Y(n3824) );
  OAI2BB2X1 U6260 ( .B0(n5515), .B1(n4931), .A0N(n5384), .A1N(x_matrix[475]), 
        .Y(n3760) );
  OAI2BB2X1 U6261 ( .B0(n5528), .B1(n4931), .A0N(n5154), .A1N(x_matrix[539]), 
        .Y(n3696) );
  OAI2BB2X1 U6262 ( .B0(n5537), .B1(n4931), .A0N(n5163), .A1N(x_matrix[587]), 
        .Y(n3632) );
  OAI2BB2X1 U6263 ( .B0(n5572), .B1(n4931), .A0N(n5171), .A1N(x_matrix[699]), 
        .Y(n3504) );
  OAI2BB2X1 U6264 ( .B0(n5407), .B1(n4929), .A0N(n5092), .A1N(x_matrix[60]), 
        .Y(n4399) );
  OAI2BB2X1 U6265 ( .B0(n5429), .B1(n4929), .A0N(n5102), .A1N(x_matrix[140]), 
        .Y(n4271) );
  OAI2BB2X1 U6266 ( .B0(n5461), .B1(n4929), .A0N(n5119), .A1N(x_matrix[252]), 
        .Y(n4079) );
  OAI2BB2X1 U6267 ( .B0(n5483), .B1(n4929), .A0N(n5135), .A1N(x_matrix[348]), 
        .Y(n3951) );
  OAI2BB2X1 U6268 ( .B0(n5494), .B1(n4929), .A0N(n5362), .A1N(x_matrix[380]), 
        .Y(n3887) );
  OAI2BB2X1 U6269 ( .B0(n5506), .B1(n4929), .A0N(n5144), .A1N(x_matrix[444]), 
        .Y(n3823) );
  OAI2BB2X1 U6270 ( .B0(n5516), .B1(n4929), .A0N(n5384), .A1N(x_matrix[476]), 
        .Y(n3759) );
  OAI2BB2X1 U6271 ( .B0(n5529), .B1(n4929), .A0N(n5155), .A1N(x_matrix[540]), 
        .Y(n3695) );
  OAI2BB2X1 U6272 ( .B0(n5538), .B1(n4929), .A0N(n5163), .A1N(x_matrix[588]), 
        .Y(n3631) );
  OAI2BB2X1 U6273 ( .B0(n5573), .B1(n4929), .A0N(n5171), .A1N(x_matrix[700]), 
        .Y(n3503) );
  OAI2BB2X1 U6274 ( .B0(n5407), .B1(n4928), .A0N(n5092), .A1N(x_matrix[61]), 
        .Y(n4398) );
  OAI2BB2X1 U6275 ( .B0(n5429), .B1(n4928), .A0N(n5102), .A1N(x_matrix[141]), 
        .Y(n4270) );
  OAI2BB2X1 U6276 ( .B0(n5460), .B1(n4928), .A0N(n5119), .A1N(x_matrix[253]), 
        .Y(n4078) );
  OAI2BB2X1 U6277 ( .B0(n5482), .B1(n4928), .A0N(n5135), .A1N(x_matrix[349]), 
        .Y(n3950) );
  OAI2BB2X1 U6278 ( .B0(n5493), .B1(n4928), .A0N(n5362), .A1N(x_matrix[381]), 
        .Y(n3886) );
  OAI2BB2X1 U6279 ( .B0(n5506), .B1(n4928), .A0N(n5144), .A1N(x_matrix[445]), 
        .Y(n3822) );
  OAI2BB2X1 U6280 ( .B0(n5515), .B1(n4928), .A0N(n5384), .A1N(x_matrix[477]), 
        .Y(n3758) );
  OAI2BB2X1 U6281 ( .B0(n5529), .B1(n4928), .A0N(n5155), .A1N(x_matrix[541]), 
        .Y(n3694) );
  OAI2BB2X1 U6282 ( .B0(n5537), .B1(n4928), .A0N(n5163), .A1N(x_matrix[589]), 
        .Y(n3630) );
  OAI2BB2X1 U6283 ( .B0(n5572), .B1(n4928), .A0N(n5171), .A1N(x_matrix[701]), 
        .Y(n3502) );
  OAI2BB2X1 U6284 ( .B0(n5407), .B1(n4927), .A0N(n5092), .A1N(x_matrix[62]), 
        .Y(n4397) );
  OAI2BB2X1 U6285 ( .B0(n5429), .B1(n4927), .A0N(n5102), .A1N(x_matrix[142]), 
        .Y(n4269) );
  OAI2BB2X1 U6286 ( .B0(n5461), .B1(n4927), .A0N(n5119), .A1N(x_matrix[254]), 
        .Y(n4077) );
  OAI2BB2X1 U6287 ( .B0(n5483), .B1(n4927), .A0N(n5135), .A1N(x_matrix[350]), 
        .Y(n3949) );
  OAI2BB2X1 U6288 ( .B0(n5493), .B1(n4927), .A0N(n5362), .A1N(x_matrix[382]), 
        .Y(n3885) );
  OAI2BB2X1 U6289 ( .B0(n5506), .B1(n4927), .A0N(n5144), .A1N(x_matrix[446]), 
        .Y(n3821) );
  OAI2BB2X1 U6290 ( .B0(n5515), .B1(n4927), .A0N(n5384), .A1N(x_matrix[478]), 
        .Y(n3757) );
  OAI2BB2X1 U6291 ( .B0(n5529), .B1(n4927), .A0N(n5155), .A1N(x_matrix[542]), 
        .Y(n3693) );
  OAI2BB2X1 U6292 ( .B0(n5538), .B1(n4927), .A0N(n5163), .A1N(x_matrix[590]), 
        .Y(n3629) );
  OAI2BB2X1 U6293 ( .B0(n5573), .B1(n4927), .A0N(n5171), .A1N(x_matrix[702]), 
        .Y(n3501) );
  OAI2BB2X1 U6294 ( .B0(n5407), .B1(n4926), .A0N(n5092), .A1N(x_matrix[63]), 
        .Y(n4396) );
  OAI2BB2X1 U6295 ( .B0(n5429), .B1(n4926), .A0N(n5102), .A1N(x_matrix[143]), 
        .Y(n4268) );
  OAI2BB2X1 U6296 ( .B0(n5459), .B1(n4926), .A0N(n5119), .A1N(x_matrix[255]), 
        .Y(n4076) );
  OAI2BB2X1 U6297 ( .B0(n5481), .B1(n4926), .A0N(n5135), .A1N(x_matrix[351]), 
        .Y(n3948) );
  OAI2BB2X1 U6298 ( .B0(n5493), .B1(n4926), .A0N(n5362), .A1N(x_matrix[383]), 
        .Y(n3884) );
  OAI2BB2X1 U6299 ( .B0(n5506), .B1(n4926), .A0N(n5144), .A1N(x_matrix[447]), 
        .Y(n3820) );
  OAI2BB2X1 U6300 ( .B0(n5515), .B1(n4926), .A0N(n5384), .A1N(x_matrix[479]), 
        .Y(n3756) );
  OAI2BB2X1 U6301 ( .B0(n5529), .B1(n4926), .A0N(n5155), .A1N(x_matrix[543]), 
        .Y(n3692) );
  OAI2BB2X1 U6302 ( .B0(n5536), .B1(n4926), .A0N(n5163), .A1N(x_matrix[591]), 
        .Y(n3628) );
  OAI2BB2X1 U6303 ( .B0(n5571), .B1(n4926), .A0N(n5171), .A1N(x_matrix[703]), 
        .Y(n3500) );
  OAI2BB2X1 U6304 ( .B0(n5405), .B1(n4960), .A0N(n5090), .A1N(x_matrix[32]), 
        .Y(n4427) );
  OAI2BB2X1 U6305 ( .B0(n5427), .B1(n4960), .A0N(n5100), .A1N(x_matrix[112]), 
        .Y(n4299) );
  OAI2BB2X1 U6306 ( .B0(n5453), .B1(n4960), .A0N(n5111), .A1N(x_matrix[192]), 
        .Y(n4171) );
  OAI2BB2X1 U6307 ( .B0(n5459), .B1(n4960), .A0N(n5118), .A1N(x_matrix[224]), 
        .Y(n4107) );
  OAI2BB2X1 U6308 ( .B0(n5475), .B1(n4960), .A0N(n5127), .A1N(x_matrix[288]), 
        .Y(n4043) );
  OAI2BB2X1 U6309 ( .B0(n5481), .B1(n4960), .A0N(n5133), .A1N(x_matrix[320]), 
        .Y(n3979) );
  OAI2BB2X1 U6310 ( .B0(n5504), .B1(n4960), .A0N(n5142), .A1N(x_matrix[416]), 
        .Y(n3851) );
  OAI2BB2X1 U6311 ( .B0(n5526), .B1(n4960), .A0N(n5153), .A1N(x_matrix[512]), 
        .Y(n3723) );
  OAI2BB2X1 U6312 ( .B0(n5536), .B1(n4960), .A0N(n5162), .A1N(x_matrix[560]), 
        .Y(n3659) );
  OAI2BB2X1 U6313 ( .B0(n5571), .B1(n4960), .A0N(n5170), .A1N(x_matrix[672]), 
        .Y(n3531) );
  OAI2BB2X1 U6314 ( .B0(n5406), .B1(n4959), .A0N(n5090), .A1N(x_matrix[33]), 
        .Y(n4426) );
  OAI2BB2X1 U6315 ( .B0(n5428), .B1(n4959), .A0N(n5100), .A1N(x_matrix[113]), 
        .Y(n4298) );
  OAI2BB2X1 U6316 ( .B0(n5452), .B1(n4959), .A0N(n5111), .A1N(x_matrix[193]), 
        .Y(n4170) );
  OAI2BB2X1 U6317 ( .B0(n5459), .B1(n4959), .A0N(n5118), .A1N(x_matrix[225]), 
        .Y(n4106) );
  OAI2BB2X1 U6318 ( .B0(n5474), .B1(n4959), .A0N(n5127), .A1N(x_matrix[289]), 
        .Y(n4042) );
  OAI2BB2X1 U6319 ( .B0(n5481), .B1(n4959), .A0N(n5133), .A1N(x_matrix[321]), 
        .Y(n3978) );
  OAI2BB2X1 U6320 ( .B0(n5505), .B1(n4959), .A0N(n5142), .A1N(x_matrix[417]), 
        .Y(n3850) );
  OAI2BB2X1 U6321 ( .B0(n5526), .B1(n4959), .A0N(n5153), .A1N(x_matrix[513]), 
        .Y(n3722) );
  OAI2BB2X1 U6322 ( .B0(n5536), .B1(n4959), .A0N(n5162), .A1N(x_matrix[561]), 
        .Y(n3658) );
  OAI2BB2X1 U6323 ( .B0(n5571), .B1(n4959), .A0N(n5170), .A1N(x_matrix[673]), 
        .Y(n3530) );
  OAI2BB2X1 U6324 ( .B0(n5405), .B1(n4958), .A0N(n5090), .A1N(x_matrix[34]), 
        .Y(n4425) );
  OAI2BB2X1 U6325 ( .B0(n5427), .B1(n4958), .A0N(n5100), .A1N(x_matrix[114]), 
        .Y(n4297) );
  OAI2BB2X1 U6326 ( .B0(n5451), .B1(n4958), .A0N(n5111), .A1N(x_matrix[194]), 
        .Y(n4169) );
  OAI2BB2X1 U6327 ( .B0(n5459), .B1(n4958), .A0N(n5118), .A1N(x_matrix[226]), 
        .Y(n4105) );
  OAI2BB2X1 U6328 ( .B0(n5473), .B1(n4958), .A0N(n5127), .A1N(x_matrix[290]), 
        .Y(n4041) );
  OAI2BB2X1 U6329 ( .B0(n5481), .B1(n4958), .A0N(n5133), .A1N(x_matrix[322]), 
        .Y(n3977) );
  OAI2BB2X1 U6330 ( .B0(n5504), .B1(n4958), .A0N(n5142), .A1N(x_matrix[418]), 
        .Y(n3849) );
  OAI2BB2X1 U6331 ( .B0(n5526), .B1(n4958), .A0N(n5153), .A1N(x_matrix[514]), 
        .Y(n3721) );
  OAI2BB2X1 U6332 ( .B0(n5536), .B1(n4958), .A0N(n5162), .A1N(x_matrix[562]), 
        .Y(n3657) );
  OAI2BB2X1 U6333 ( .B0(n5571), .B1(n4958), .A0N(n5170), .A1N(x_matrix[674]), 
        .Y(n3529) );
  OAI2BB2X1 U6334 ( .B0(n5406), .B1(n4957), .A0N(n5090), .A1N(x_matrix[35]), 
        .Y(n4424) );
  OAI2BB2X1 U6335 ( .B0(n5428), .B1(n4957), .A0N(n5100), .A1N(x_matrix[115]), 
        .Y(n4296) );
  OAI2BB2X1 U6336 ( .B0(n5453), .B1(n4957), .A0N(n5111), .A1N(x_matrix[195]), 
        .Y(n4168) );
  OAI2BB2X1 U6337 ( .B0(n5459), .B1(n4957), .A0N(n5118), .A1N(x_matrix[227]), 
        .Y(n4104) );
  OAI2BB2X1 U6338 ( .B0(n5475), .B1(n4957), .A0N(n5127), .A1N(x_matrix[291]), 
        .Y(n4040) );
  OAI2BB2X1 U6339 ( .B0(n5481), .B1(n4957), .A0N(n5133), .A1N(x_matrix[323]), 
        .Y(n3976) );
  OAI2BB2X1 U6340 ( .B0(n5505), .B1(n4957), .A0N(n5142), .A1N(x_matrix[419]), 
        .Y(n3848) );
  OAI2BB2X1 U6341 ( .B0(n5526), .B1(n4957), .A0N(n5153), .A1N(x_matrix[515]), 
        .Y(n3720) );
  OAI2BB2X1 U6342 ( .B0(n5536), .B1(n4957), .A0N(n5162), .A1N(x_matrix[563]), 
        .Y(n3656) );
  OAI2BB2X1 U6343 ( .B0(n5571), .B1(n4957), .A0N(n5170), .A1N(x_matrix[675]), 
        .Y(n3528) );
  OAI2BB2X1 U6344 ( .B0(n5405), .B1(n4956), .A0N(n5091), .A1N(x_matrix[36]), 
        .Y(n4423) );
  OAI2BB2X1 U6345 ( .B0(n5427), .B1(n4956), .A0N(n5101), .A1N(x_matrix[116]), 
        .Y(n4295) );
  OAI2BB2X1 U6346 ( .B0(n5450), .B1(n4956), .A0N(n5111), .A1N(x_matrix[196]), 
        .Y(n4167) );
  OAI2BB2X1 U6347 ( .B0(n5459), .B1(n4956), .A0N(n5118), .A1N(x_matrix[228]), 
        .Y(n4103) );
  OAI2BB2X1 U6348 ( .B0(n5472), .B1(n4956), .A0N(n5127), .A1N(x_matrix[292]), 
        .Y(n4039) );
  OAI2BB2X1 U6349 ( .B0(n5481), .B1(n4956), .A0N(n5133), .A1N(x_matrix[324]), 
        .Y(n3975) );
  OAI2BB2X1 U6350 ( .B0(n5504), .B1(n4956), .A0N(n5143), .A1N(x_matrix[420]), 
        .Y(n3847) );
  OAI2BB2X1 U6351 ( .B0(n5527), .B1(n4956), .A0N(n5152), .A1N(x_matrix[516]), 
        .Y(n3719) );
  OAI2BB2X1 U6352 ( .B0(n5536), .B1(n4956), .A0N(n5162), .A1N(x_matrix[564]), 
        .Y(n3655) );
  OAI2BB2X1 U6353 ( .B0(n5571), .B1(n4956), .A0N(n5170), .A1N(x_matrix[676]), 
        .Y(n3527) );
  OAI2BB2X1 U6354 ( .B0(n5405), .B1(n4955), .A0N(n5091), .A1N(x_matrix[37]), 
        .Y(n4422) );
  OAI2BB2X1 U6355 ( .B0(n5427), .B1(n4955), .A0N(n5101), .A1N(x_matrix[117]), 
        .Y(n4294) );
  OAI2BB2X1 U6356 ( .B0(n5450), .B1(n4955), .A0N(n5111), .A1N(x_matrix[197]), 
        .Y(n4166) );
  OAI2BB2X1 U6357 ( .B0(n5459), .B1(n4955), .A0N(n5118), .A1N(x_matrix[229]), 
        .Y(n4102) );
  OAI2BB2X1 U6358 ( .B0(n5472), .B1(n4955), .A0N(n5127), .A1N(x_matrix[293]), 
        .Y(n4038) );
  OAI2BB2X1 U6359 ( .B0(n5481), .B1(n4955), .A0N(n5133), .A1N(x_matrix[325]), 
        .Y(n3974) );
  OAI2BB2X1 U6360 ( .B0(n5504), .B1(n4955), .A0N(n5143), .A1N(x_matrix[421]), 
        .Y(n3846) );
  OAI2BB2X1 U6361 ( .B0(n5527), .B1(n4955), .A0N(n5153), .A1N(x_matrix[517]), 
        .Y(n3718) );
  OAI2BB2X1 U6362 ( .B0(n5536), .B1(n4955), .A0N(n5162), .A1N(x_matrix[565]), 
        .Y(n3654) );
  OAI2BB2X1 U6363 ( .B0(n5571), .B1(n4955), .A0N(n5170), .A1N(x_matrix[677]), 
        .Y(n3526) );
  OAI2BB2X1 U6364 ( .B0(n5405), .B1(n4954), .A0N(n5091), .A1N(x_matrix[38]), 
        .Y(n4421) );
  OAI2BB2X1 U6365 ( .B0(n5427), .B1(n4954), .A0N(n5101), .A1N(x_matrix[118]), 
        .Y(n4293) );
  OAI2BB2X1 U6366 ( .B0(n5450), .B1(n4954), .A0N(n5111), .A1N(x_matrix[198]), 
        .Y(n4165) );
  OAI2BB2X1 U6367 ( .B0(n5459), .B1(n4954), .A0N(n5118), .A1N(x_matrix[230]), 
        .Y(n4101) );
  OAI2BB2X1 U6368 ( .B0(n5472), .B1(n4954), .A0N(n5127), .A1N(x_matrix[294]), 
        .Y(n4037) );
  OAI2BB2X1 U6369 ( .B0(n5481), .B1(n4954), .A0N(n5133), .A1N(x_matrix[326]), 
        .Y(n3973) );
  OAI2BB2X1 U6370 ( .B0(n5504), .B1(n4954), .A0N(n5143), .A1N(x_matrix[422]), 
        .Y(n3845) );
  OAI2BB2X1 U6371 ( .B0(n5527), .B1(n4954), .A0N(n5154), .A1N(x_matrix[518]), 
        .Y(n3717) );
  OAI2BB2X1 U6372 ( .B0(n5536), .B1(n4954), .A0N(n5162), .A1N(x_matrix[566]), 
        .Y(n3653) );
  OAI2BB2X1 U6373 ( .B0(n5571), .B1(n4954), .A0N(n5170), .A1N(x_matrix[678]), 
        .Y(n3525) );
  OAI2BB2X1 U6374 ( .B0(n5405), .B1(n4953), .A0N(n5091), .A1N(x_matrix[39]), 
        .Y(n4420) );
  OAI2BB2X1 U6375 ( .B0(n5427), .B1(n4953), .A0N(n5101), .A1N(x_matrix[119]), 
        .Y(n4292) );
  OAI2BB2X1 U6376 ( .B0(n5450), .B1(n4953), .A0N(n5111), .A1N(x_matrix[199]), 
        .Y(n4164) );
  OAI2BB2X1 U6377 ( .B0(n5459), .B1(n4953), .A0N(n5118), .A1N(x_matrix[231]), 
        .Y(n4100) );
  OAI2BB2X1 U6378 ( .B0(n5472), .B1(n4953), .A0N(n5127), .A1N(x_matrix[295]), 
        .Y(n4036) );
  OAI2BB2X1 U6379 ( .B0(n5481), .B1(n4953), .A0N(n5133), .A1N(x_matrix[327]), 
        .Y(n3972) );
  OAI2BB2X1 U6380 ( .B0(n5504), .B1(n4953), .A0N(n5143), .A1N(x_matrix[423]), 
        .Y(n3844) );
  OAI2BB2X1 U6381 ( .B0(n5527), .B1(n4953), .A0N(n5152), .A1N(x_matrix[519]), 
        .Y(n3716) );
  OAI2BB2X1 U6382 ( .B0(n5536), .B1(n4953), .A0N(n5162), .A1N(x_matrix[567]), 
        .Y(n3652) );
  OAI2BB2X1 U6383 ( .B0(n5571), .B1(n4953), .A0N(n5170), .A1N(x_matrix[679]), 
        .Y(n3524) );
  OAI2BB2X1 U6384 ( .B0(n5405), .B1(n4951), .A0N(n5091), .A1N(x_matrix[40]), 
        .Y(n4419) );
  OAI2BB2X1 U6385 ( .B0(n5427), .B1(n4951), .A0N(n5101), .A1N(x_matrix[120]), 
        .Y(n4291) );
  OAI2BB2X1 U6386 ( .B0(n5448), .B1(n4951), .A0N(n5109), .A1N(x_matrix[200]), 
        .Y(n4163) );
  OAI2BB2X1 U6387 ( .B0(n5459), .B1(n4951), .A0N(n5117), .A1N(x_matrix[232]), 
        .Y(n4099) );
  OAI2BB2X1 U6388 ( .B0(n5470), .B1(n4951), .A0N(n5125), .A1N(x_matrix[296]), 
        .Y(n4035) );
  OAI2BB2X1 U6389 ( .B0(n5481), .B1(n4951), .A0N(n5134), .A1N(x_matrix[328]), 
        .Y(n3971) );
  OAI2BB2X1 U6390 ( .B0(n5504), .B1(n4951), .A0N(n5143), .A1N(x_matrix[424]), 
        .Y(n3843) );
  OAI2BB2X1 U6391 ( .B0(n5527), .B1(n4951), .A0N(n5153), .A1N(x_matrix[520]), 
        .Y(n3715) );
  OAI2BB2X1 U6392 ( .B0(n5536), .B1(n4951), .A0N(n5161), .A1N(x_matrix[568]), 
        .Y(n3651) );
  OAI2BB2X1 U6393 ( .B0(n5571), .B1(n4951), .A0N(n5169), .A1N(x_matrix[680]), 
        .Y(n3523) );
  OAI2BB2X1 U6394 ( .B0(n5405), .B1(n4950), .A0N(n5091), .A1N(x_matrix[41]), 
        .Y(n4418) );
  OAI2BB2X1 U6395 ( .B0(n5427), .B1(n4950), .A0N(n5101), .A1N(x_matrix[121]), 
        .Y(n4290) );
  OAI2BB2X1 U6396 ( .B0(n5448), .B1(n4950), .A0N(n5110), .A1N(x_matrix[201]), 
        .Y(n4162) );
  OAI2BB2X1 U6397 ( .B0(n5465), .B1(n4950), .A0N(n5118), .A1N(x_matrix[233]), 
        .Y(n4098) );
  OAI2BB2X1 U6398 ( .B0(n5470), .B1(n4950), .A0N(n5126), .A1N(x_matrix[297]), 
        .Y(n4034) );
  OAI2BB2X1 U6399 ( .B0(n5487), .B1(n4950), .A0N(n5134), .A1N(x_matrix[329]), 
        .Y(n3970) );
  OAI2BB2X1 U6400 ( .B0(n5504), .B1(n4950), .A0N(n5143), .A1N(x_matrix[425]), 
        .Y(n3842) );
  OAI2BB2X1 U6401 ( .B0(n5527), .B1(n4950), .A0N(n5154), .A1N(x_matrix[521]), 
        .Y(n3714) );
  OAI2BB2X1 U6402 ( .B0(n5542), .B1(n4950), .A0N(n5162), .A1N(x_matrix[569]), 
        .Y(n3650) );
  OAI2BB2X1 U6403 ( .B0(n5577), .B1(n4950), .A0N(n5170), .A1N(x_matrix[681]), 
        .Y(n3522) );
  OAI2BB2X1 U6404 ( .B0(n5405), .B1(n4949), .A0N(n5091), .A1N(x_matrix[42]), 
        .Y(n4417) );
  OAI2BB2X1 U6405 ( .B0(n5427), .B1(n4949), .A0N(n5101), .A1N(x_matrix[122]), 
        .Y(n4289) );
  OAI2BB2X1 U6406 ( .B0(n5448), .B1(n4949), .A0N(n5109), .A1N(x_matrix[202]), 
        .Y(n4161) );
  OAI2BB2X1 U6407 ( .B0(n5459), .B1(n4949), .A0N(n5117), .A1N(x_matrix[234]), 
        .Y(n4097) );
  OAI2BB2X1 U6408 ( .B0(n5470), .B1(n4949), .A0N(n5125), .A1N(x_matrix[298]), 
        .Y(n4033) );
  OAI2BB2X1 U6409 ( .B0(n5481), .B1(n4949), .A0N(n5134), .A1N(x_matrix[330]), 
        .Y(n3969) );
  OAI2BB2X1 U6410 ( .B0(n5504), .B1(n4949), .A0N(n5143), .A1N(x_matrix[426]), 
        .Y(n3841) );
  OAI2BB2X1 U6411 ( .B0(n5527), .B1(n4949), .A0N(n5152), .A1N(x_matrix[522]), 
        .Y(n3713) );
  OAI2BB2X1 U6412 ( .B0(n5536), .B1(n4949), .A0N(n5161), .A1N(x_matrix[570]), 
        .Y(n3649) );
  OAI2BB2X1 U6413 ( .B0(n5571), .B1(n4949), .A0N(n5169), .A1N(x_matrix[682]), 
        .Y(n3521) );
  OAI2BB2X1 U6414 ( .B0(n5405), .B1(n4948), .A0N(n5091), .A1N(x_matrix[43]), 
        .Y(n4416) );
  OAI2BB2X1 U6415 ( .B0(n5427), .B1(n4948), .A0N(n5101), .A1N(x_matrix[123]), 
        .Y(n4288) );
  OAI2BB2X1 U6416 ( .B0(n5455), .B1(n4948), .A0N(n5110), .A1N(x_matrix[203]), 
        .Y(n4160) );
  OAI2BB2X1 U6417 ( .B0(n5465), .B1(n4948), .A0N(n5118), .A1N(x_matrix[235]), 
        .Y(n4096) );
  OAI2BB2X1 U6418 ( .B0(n5477), .B1(n4948), .A0N(n5126), .A1N(x_matrix[299]), 
        .Y(n4032) );
  OAI2BB2X1 U6419 ( .B0(n5487), .B1(n4948), .A0N(n5134), .A1N(x_matrix[331]), 
        .Y(n3968) );
  OAI2BB2X1 U6420 ( .B0(n5504), .B1(n4948), .A0N(n5143), .A1N(x_matrix[427]), 
        .Y(n3840) );
  OAI2BB2X1 U6421 ( .B0(n5527), .B1(n4948), .A0N(n5153), .A1N(x_matrix[523]), 
        .Y(n3712) );
  OAI2BB2X1 U6422 ( .B0(n5542), .B1(n4948), .A0N(n5162), .A1N(x_matrix[571]), 
        .Y(n3648) );
  OAI2BB2X1 U6423 ( .B0(n5577), .B1(n4948), .A0N(n5170), .A1N(x_matrix[683]), 
        .Y(n3520) );
  OAI2BB2X1 U6424 ( .B0(n5405), .B1(n4947), .A0N(n5091), .A1N(x_matrix[44]), 
        .Y(n4415) );
  OAI2BB2X1 U6425 ( .B0(n5427), .B1(n4947), .A0N(n5101), .A1N(x_matrix[124]), 
        .Y(n4287) );
  OAI2BB2X1 U6426 ( .B0(n5448), .B1(n4947), .A0N(n5109), .A1N(x_matrix[204]), 
        .Y(n4159) );
  OAI2BB2X1 U6427 ( .B0(n5464), .B1(n4947), .A0N(n5117), .A1N(x_matrix[236]), 
        .Y(n4095) );
  OAI2BB2X1 U6428 ( .B0(n5470), .B1(n4947), .A0N(n5125), .A1N(x_matrix[300]), 
        .Y(n4031) );
  OAI2BB2X1 U6429 ( .B0(n5486), .B1(n4947), .A0N(n5134), .A1N(x_matrix[332]), 
        .Y(n3967) );
  OAI2BB2X1 U6430 ( .B0(n5504), .B1(n4947), .A0N(n5143), .A1N(x_matrix[428]), 
        .Y(n3839) );
  OAI2BB2X1 U6431 ( .B0(n5527), .B1(n4947), .A0N(n5154), .A1N(x_matrix[524]), 
        .Y(n3711) );
  OAI2BB2X1 U6432 ( .B0(n5541), .B1(n4947), .A0N(n5161), .A1N(x_matrix[572]), 
        .Y(n3647) );
  OAI2BB2X1 U6433 ( .B0(n5576), .B1(n4947), .A0N(n5169), .A1N(x_matrix[684]), 
        .Y(n3519) );
  OAI2BB2X1 U6434 ( .B0(n5405), .B1(n4946), .A0N(n5091), .A1N(x_matrix[45]), 
        .Y(n4414) );
  OAI2BB2X1 U6435 ( .B0(n5427), .B1(n4946), .A0N(n5101), .A1N(x_matrix[125]), 
        .Y(n4286) );
  OAI2BB2X1 U6436 ( .B0(n5455), .B1(n4946), .A0N(n5110), .A1N(x_matrix[205]), 
        .Y(n4158) );
  OAI2BB2X1 U6437 ( .B0(n5463), .B1(n4946), .A0N(n5118), .A1N(x_matrix[237]), 
        .Y(n4094) );
  OAI2BB2X1 U6438 ( .B0(n5477), .B1(n4946), .A0N(n5126), .A1N(x_matrix[301]), 
        .Y(n4030) );
  OAI2BB2X1 U6439 ( .B0(n5485), .B1(n4946), .A0N(n5134), .A1N(x_matrix[333]), 
        .Y(n3966) );
  OAI2BB2X1 U6440 ( .B0(n5504), .B1(n4946), .A0N(n5143), .A1N(x_matrix[429]), 
        .Y(n3838) );
  OAI2BB2X1 U6441 ( .B0(n5527), .B1(n4946), .A0N(n5152), .A1N(x_matrix[525]), 
        .Y(n3710) );
  OAI2BB2X1 U6442 ( .B0(n5540), .B1(n4946), .A0N(n5162), .A1N(x_matrix[573]), 
        .Y(n3646) );
  OAI2BB2X1 U6443 ( .B0(n5575), .B1(n4946), .A0N(n5170), .A1N(x_matrix[685]), 
        .Y(n3518) );
  OAI2BB2X1 U6444 ( .B0(n5405), .B1(n4945), .A0N(n5091), .A1N(x_matrix[46]), 
        .Y(n4413) );
  OAI2BB2X1 U6445 ( .B0(n5427), .B1(n4945), .A0N(n5101), .A1N(x_matrix[126]), 
        .Y(n4285) );
  OAI2BB2X1 U6446 ( .B0(n5448), .B1(n4945), .A0N(n5116), .A1N(x_matrix[206]), 
        .Y(n4157) );
  OAI2BB2X1 U6447 ( .B0(n5462), .B1(n4945), .A0N(n5124), .A1N(x_matrix[238]), 
        .Y(n4093) );
  OAI2BB2X1 U6448 ( .B0(n5470), .B1(n4945), .A0N(n5132), .A1N(x_matrix[302]), 
        .Y(n4029) );
  OAI2BB2X1 U6449 ( .B0(n5484), .B1(n4945), .A0N(n5134), .A1N(x_matrix[334]), 
        .Y(n3965) );
  OAI2BB2X1 U6450 ( .B0(n5504), .B1(n4945), .A0N(n5143), .A1N(x_matrix[430]), 
        .Y(n3837) );
  OAI2BB2X1 U6451 ( .B0(n5527), .B1(n4945), .A0N(n5153), .A1N(x_matrix[526]), 
        .Y(n3709) );
  OAI2BB2X1 U6452 ( .B0(n5539), .B1(n4945), .A0N(n5168), .A1N(x_matrix[574]), 
        .Y(n3645) );
  OAI2BB2X1 U6453 ( .B0(n5574), .B1(n4945), .A0N(n5176), .A1N(x_matrix[686]), 
        .Y(n3517) );
  OAI2BB2X1 U6454 ( .B0(n5405), .B1(n4944), .A0N(n5091), .A1N(x_matrix[47]), 
        .Y(n4412) );
  OAI2BB2X1 U6455 ( .B0(n5427), .B1(n4944), .A0N(n5101), .A1N(x_matrix[127]), 
        .Y(n4284) );
  OAI2BB2X1 U6456 ( .B0(n5449), .B1(n4944), .A0N(n5109), .A1N(x_matrix[207]), 
        .Y(n4156) );
  OAI2BB2X1 U6457 ( .B0(n5464), .B1(n4944), .A0N(n5117), .A1N(x_matrix[239]), 
        .Y(n4092) );
  OAI2BB2X1 U6458 ( .B0(n5471), .B1(n4944), .A0N(n5125), .A1N(x_matrix[303]), 
        .Y(n4028) );
  OAI2BB2X1 U6459 ( .B0(n5486), .B1(n4944), .A0N(n5134), .A1N(x_matrix[335]), 
        .Y(n3964) );
  OAI2BB2X1 U6460 ( .B0(n5504), .B1(n4944), .A0N(n5143), .A1N(x_matrix[431]), 
        .Y(n3836) );
  OAI2BB2X1 U6461 ( .B0(n5527), .B1(n4944), .A0N(n5154), .A1N(x_matrix[527]), 
        .Y(n3708) );
  OAI2BB2X1 U6462 ( .B0(n5541), .B1(n4944), .A0N(n5161), .A1N(x_matrix[575]), 
        .Y(n3644) );
  OAI2BB2X1 U6463 ( .B0(n5576), .B1(n4944), .A0N(n5169), .A1N(x_matrix[687]), 
        .Y(n3516) );
  OAI2BB2X1 U6464 ( .B0(n5049), .B1(n5461), .A0N(w_matrix[320]), .A1N(n5120), 
        .Y(n3115) );
  OAI2BB2X1 U6465 ( .B0(n5049), .B1(n5483), .A0N(w_matrix[448]), .A1N(n5136), 
        .Y(n2987) );
  OAI2BB2X1 U6466 ( .B0(n5049), .B1(n5538), .A0N(w_matrix[768]), .A1N(n5164), 
        .Y(n2667) );
  OAI2BB2X1 U6467 ( .B0(n5049), .B1(n5573), .A0N(w_matrix[896]), .A1N(n5172), 
        .Y(n2539) );
  OAI2BB2X1 U6468 ( .B0(n5048), .B1(n5408), .A0N(w_matrix[10]), .A1N(n5093), 
        .Y(n3425) );
  OAI2BB2X1 U6469 ( .B0(n5048), .B1(n5430), .A0N(w_matrix[138]), .A1N(n5103), 
        .Y(n3297) );
  OAI2BB2X1 U6470 ( .B0(n5048), .B1(n5462), .A0N(w_matrix[330]), .A1N(n5120), 
        .Y(n3105) );
  OAI2BB2X1 U6471 ( .B0(n5048), .B1(n5484), .A0N(w_matrix[458]), .A1N(n5136), 
        .Y(n2977) );
  OAI2BB2X1 U6472 ( .B0(n5048), .B1(n5507), .A0N(w_matrix[586]), .A1N(n5145), 
        .Y(n2849) );
  OAI2BB2X1 U6473 ( .B0(n5048), .B1(n5529), .A0N(w_matrix[714]), .A1N(n5156), 
        .Y(n2721) );
  OAI2BB2X1 U6474 ( .B0(n5048), .B1(n5539), .A0N(w_matrix[778]), .A1N(n5164), 
        .Y(n2657) );
  OAI2BB2X1 U6475 ( .B0(n5048), .B1(n5574), .A0N(w_matrix[906]), .A1N(n5172), 
        .Y(n2529) );
  OAI2BB2X1 U6476 ( .B0(n5047), .B1(n5408), .A0N(w_matrix[11]), .A1N(n5093), 
        .Y(n3424) );
  OAI2BB2X1 U6477 ( .B0(n5047), .B1(n5430), .A0N(w_matrix[139]), .A1N(n5103), 
        .Y(n3296) );
  OAI2BB2X1 U6478 ( .B0(n5047), .B1(n5462), .A0N(w_matrix[331]), .A1N(n5120), 
        .Y(n3104) );
  OAI2BB2X1 U6479 ( .B0(n5047), .B1(n5484), .A0N(w_matrix[459]), .A1N(n5136), 
        .Y(n2976) );
  OAI2BB2X1 U6480 ( .B0(n5047), .B1(n5507), .A0N(w_matrix[587]), .A1N(n5145), 
        .Y(n2848) );
  OAI2BB2X1 U6481 ( .B0(n5047), .B1(n5531), .A0N(w_matrix[715]), .A1N(n5156), 
        .Y(n2720) );
  OAI2BB2X1 U6482 ( .B0(n5047), .B1(n5539), .A0N(w_matrix[779]), .A1N(n5164), 
        .Y(n2656) );
  OAI2BB2X1 U6483 ( .B0(n5047), .B1(n5574), .A0N(w_matrix[907]), .A1N(n5172), 
        .Y(n2528) );
  OAI2BB2X1 U6484 ( .B0(n5046), .B1(n5408), .A0N(w_matrix[12]), .A1N(n5093), 
        .Y(n3423) );
  OAI2BB2X1 U6485 ( .B0(n5046), .B1(n5430), .A0N(w_matrix[140]), .A1N(n5103), 
        .Y(n3295) );
  OAI2BB2X1 U6486 ( .B0(n5046), .B1(n5453), .A0N(w_matrix[268]), .A1N(n5112), 
        .Y(n3167) );
  OAI2BB2X1 U6487 ( .B0(n5046), .B1(n5461), .A0N(w_matrix[332]), .A1N(n5120), 
        .Y(n3103) );
  OAI2BB2X1 U6488 ( .B0(n5046), .B1(n5475), .A0N(w_matrix[396]), .A1N(n5128), 
        .Y(n3039) );
  OAI2BB2X1 U6489 ( .B0(n5046), .B1(n5483), .A0N(w_matrix[460]), .A1N(n5136), 
        .Y(n2975) );
  OAI2BB2X1 U6490 ( .B0(n5046), .B1(n5507), .A0N(w_matrix[588]), .A1N(n5145), 
        .Y(n2847) );
  OAI2BB2X1 U6491 ( .B0(n5046), .B1(n5529), .A0N(w_matrix[716]), .A1N(n5156), 
        .Y(n2719) );
  OAI2BB2X1 U6492 ( .B0(n5046), .B1(n5538), .A0N(w_matrix[780]), .A1N(n5164), 
        .Y(n2655) );
  OAI2BB2X1 U6493 ( .B0(n5046), .B1(n5573), .A0N(w_matrix[908]), .A1N(n5172), 
        .Y(n2527) );
  OAI2BB2X1 U6494 ( .B0(n5045), .B1(n5408), .A0N(w_matrix[13]), .A1N(n5093), 
        .Y(n3422) );
  OAI2BB2X1 U6495 ( .B0(n5045), .B1(n5430), .A0N(w_matrix[141]), .A1N(n5103), 
        .Y(n3294) );
  OAI2BB2X1 U6496 ( .B0(n5045), .B1(n5453), .A0N(w_matrix[269]), .A1N(n5113), 
        .Y(n3166) );
  OAI2BB2X1 U6497 ( .B0(n5045), .B1(n5462), .A0N(w_matrix[333]), .A1N(n5121), 
        .Y(n3102) );
  OAI2BB2X1 U6498 ( .B0(n5045), .B1(n5475), .A0N(w_matrix[397]), .A1N(n5129), 
        .Y(n3038) );
  OAI2BB2X1 U6499 ( .B0(n5045), .B1(n5484), .A0N(w_matrix[461]), .A1N(n5137), 
        .Y(n2974) );
  OAI2BB2X1 U6500 ( .B0(n5045), .B1(n5507), .A0N(w_matrix[589]), .A1N(n5145), 
        .Y(n2846) );
  OAI2BB2X1 U6501 ( .B0(n5045), .B1(n5531), .A0N(w_matrix[717]), .A1N(n5156), 
        .Y(n2718) );
  OAI2BB2X1 U6502 ( .B0(n5045), .B1(n5539), .A0N(w_matrix[781]), .A1N(n5165), 
        .Y(n2654) );
  OAI2BB2X1 U6503 ( .B0(n5045), .B1(n5574), .A0N(w_matrix[909]), .A1N(n5173), 
        .Y(n2526) );
  OAI2BB2X1 U6504 ( .B0(n5044), .B1(n5408), .A0N(w_matrix[14]), .A1N(n5093), 
        .Y(n3421) );
  OAI2BB2X1 U6505 ( .B0(n5044), .B1(n5430), .A0N(w_matrix[142]), .A1N(n5103), 
        .Y(n3293) );
  OAI2BB2X1 U6506 ( .B0(n5044), .B1(n5453), .A0N(w_matrix[270]), .A1N(n5113), 
        .Y(n3165) );
  OAI2BB2X1 U6507 ( .B0(n5044), .B1(n5462), .A0N(w_matrix[334]), .A1N(n5121), 
        .Y(n3101) );
  OAI2BB2X1 U6508 ( .B0(n5044), .B1(n5475), .A0N(w_matrix[398]), .A1N(n5129), 
        .Y(n3037) );
  OAI2BB2X1 U6509 ( .B0(n5044), .B1(n5484), .A0N(w_matrix[462]), .A1N(n5137), 
        .Y(n2973) );
  OAI2BB2X1 U6510 ( .B0(n5044), .B1(n5507), .A0N(w_matrix[590]), .A1N(n5145), 
        .Y(n2845) );
  OAI2BB2X1 U6511 ( .B0(n5044), .B1(n5529), .A0N(w_matrix[718]), .A1N(n5156), 
        .Y(n2717) );
  OAI2BB2X1 U6512 ( .B0(n5044), .B1(n5539), .A0N(w_matrix[782]), .A1N(n5165), 
        .Y(n2653) );
  OAI2BB2X1 U6513 ( .B0(n5044), .B1(n5574), .A0N(w_matrix[910]), .A1N(n5173), 
        .Y(n2525) );
  OAI2BB2X1 U6514 ( .B0(n5043), .B1(n5408), .A0N(w_matrix[15]), .A1N(n5093), 
        .Y(n3420) );
  OAI2BB2X1 U6515 ( .B0(n5043), .B1(n5430), .A0N(w_matrix[143]), .A1N(n5103), 
        .Y(n3292) );
  OAI2BB2X1 U6516 ( .B0(n5043), .B1(n5453), .A0N(w_matrix[271]), .A1N(n5113), 
        .Y(n3164) );
  OAI2BB2X1 U6517 ( .B0(n5043), .B1(n5461), .A0N(w_matrix[335]), .A1N(n5121), 
        .Y(n3100) );
  OAI2BB2X1 U6518 ( .B0(n5043), .B1(n5475), .A0N(w_matrix[399]), .A1N(n5129), 
        .Y(n3036) );
  OAI2BB2X1 U6519 ( .B0(n5043), .B1(n5483), .A0N(w_matrix[463]), .A1N(n5137), 
        .Y(n2972) );
  OAI2BB2X1 U6520 ( .B0(n5043), .B1(n5507), .A0N(w_matrix[591]), .A1N(n5145), 
        .Y(n2844) );
  OAI2BB2X1 U6521 ( .B0(n5043), .B1(n5530), .A0N(w_matrix[719]), .A1N(n5156), 
        .Y(n2716) );
  OAI2BB2X1 U6522 ( .B0(n5043), .B1(n5538), .A0N(w_matrix[783]), .A1N(n5165), 
        .Y(n2652) );
  OAI2BB2X1 U6523 ( .B0(n5043), .B1(n5573), .A0N(w_matrix[911]), .A1N(n5173), 
        .Y(n2524) );
  OAI2BB2X1 U6524 ( .B0(n5042), .B1(n5408), .A0N(w_matrix[16]), .A1N(n5093), 
        .Y(n3419) );
  OAI2BB2X1 U6525 ( .B0(n5042), .B1(n5430), .A0N(w_matrix[144]), .A1N(n5103), 
        .Y(n3291) );
  OAI2BB2X1 U6526 ( .B0(n5042), .B1(n5453), .A0N(w_matrix[272]), .A1N(n5113), 
        .Y(n3163) );
  OAI2BB2X1 U6527 ( .B0(n5042), .B1(n5462), .A0N(w_matrix[336]), .A1N(n5121), 
        .Y(n3099) );
  OAI2BB2X1 U6528 ( .B0(n5042), .B1(n5475), .A0N(w_matrix[400]), .A1N(n5129), 
        .Y(n3035) );
  OAI2BB2X1 U6529 ( .B0(n5042), .B1(n5484), .A0N(w_matrix[464]), .A1N(n5137), 
        .Y(n2971) );
  OAI2BB2X1 U6530 ( .B0(n5042), .B1(n5507), .A0N(w_matrix[592]), .A1N(n5145), 
        .Y(n2843) );
  OAI2BB2X1 U6531 ( .B0(n5042), .B1(n5525), .A0N(w_matrix[720]), .A1N(n5156), 
        .Y(n2715) );
  OAI2BB2X1 U6532 ( .B0(n5042), .B1(n5539), .A0N(w_matrix[784]), .A1N(n5165), 
        .Y(n2651) );
  OAI2BB2X1 U6533 ( .B0(n5042), .B1(n5574), .A0N(w_matrix[912]), .A1N(n5173), 
        .Y(n2523) );
  OAI2BB2X1 U6534 ( .B0(n5041), .B1(n5408), .A0N(w_matrix[17]), .A1N(n5093), 
        .Y(n3418) );
  OAI2BB2X1 U6535 ( .B0(n5041), .B1(n5430), .A0N(w_matrix[145]), .A1N(n5103), 
        .Y(n3290) );
  OAI2BB2X1 U6536 ( .B0(n5041), .B1(n5453), .A0N(w_matrix[273]), .A1N(n5113), 
        .Y(n3162) );
  OAI2BB2X1 U6537 ( .B0(n5041), .B1(n5462), .A0N(w_matrix[337]), .A1N(n5121), 
        .Y(n3098) );
  OAI2BB2X1 U6538 ( .B0(n5041), .B1(n5475), .A0N(w_matrix[401]), .A1N(n5129), 
        .Y(n3034) );
  OAI2BB2X1 U6539 ( .B0(n5041), .B1(n5484), .A0N(w_matrix[465]), .A1N(n5137), 
        .Y(n2970) );
  OAI2BB2X1 U6540 ( .B0(n5041), .B1(n5507), .A0N(w_matrix[593]), .A1N(n5145), 
        .Y(n2842) );
  OAI2BB2X1 U6541 ( .B0(n5041), .B1(n5526), .A0N(w_matrix[721]), .A1N(n5156), 
        .Y(n2714) );
  OAI2BB2X1 U6542 ( .B0(n5041), .B1(n5539), .A0N(w_matrix[785]), .A1N(n5165), 
        .Y(n2650) );
  OAI2BB2X1 U6543 ( .B0(n5041), .B1(n5574), .A0N(w_matrix[913]), .A1N(n5173), 
        .Y(n2522) );
  OAI2BB2X1 U6544 ( .B0(n5040), .B1(n5408), .A0N(w_matrix[18]), .A1N(n5093), 
        .Y(n3417) );
  OAI2BB2X1 U6545 ( .B0(n5040), .B1(n5430), .A0N(w_matrix[146]), .A1N(n5103), 
        .Y(n3289) );
  OAI2BB2X1 U6546 ( .B0(n5040), .B1(n5453), .A0N(w_matrix[274]), .A1N(n5113), 
        .Y(n3161) );
  OAI2BB2X1 U6547 ( .B0(n5040), .B1(n5462), .A0N(w_matrix[338]), .A1N(n5121), 
        .Y(n3097) );
  OAI2BB2X1 U6548 ( .B0(n5040), .B1(n5475), .A0N(w_matrix[402]), .A1N(n5129), 
        .Y(n3033) );
  OAI2BB2X1 U6549 ( .B0(n5040), .B1(n5484), .A0N(w_matrix[466]), .A1N(n5137), 
        .Y(n2969) );
  OAI2BB2X1 U6550 ( .B0(n5040), .B1(n5507), .A0N(w_matrix[594]), .A1N(n5145), 
        .Y(n2841) );
  OAI2BB2X1 U6551 ( .B0(n5040), .B1(n5527), .A0N(w_matrix[722]), .A1N(n5156), 
        .Y(n2713) );
  OAI2BB2X1 U6552 ( .B0(n5040), .B1(n5539), .A0N(w_matrix[786]), .A1N(n5165), 
        .Y(n2649) );
  OAI2BB2X1 U6553 ( .B0(n5040), .B1(n5574), .A0N(w_matrix[914]), .A1N(n5173), 
        .Y(n2521) );
  OAI2BB2X1 U6554 ( .B0(n5039), .B1(n5408), .A0N(w_matrix[19]), .A1N(n5093), 
        .Y(n3416) );
  OAI2BB2X1 U6555 ( .B0(n5039), .B1(n5430), .A0N(w_matrix[147]), .A1N(n5103), 
        .Y(n3288) );
  OAI2BB2X1 U6556 ( .B0(n5039), .B1(n5453), .A0N(w_matrix[275]), .A1N(n5113), 
        .Y(n3160) );
  OAI2BB2X1 U6557 ( .B0(n5039), .B1(n5463), .A0N(w_matrix[339]), .A1N(n5121), 
        .Y(n3096) );
  OAI2BB2X1 U6558 ( .B0(n5039), .B1(n5475), .A0N(w_matrix[403]), .A1N(n5129), 
        .Y(n3032) );
  OAI2BB2X1 U6559 ( .B0(n5039), .B1(n5485), .A0N(w_matrix[467]), .A1N(n5137), 
        .Y(n2968) );
  OAI2BB2X1 U6560 ( .B0(n5039), .B1(n5507), .A0N(w_matrix[595]), .A1N(n5145), 
        .Y(n2840) );
  OAI2BB2X1 U6561 ( .B0(n5039), .B1(n5528), .A0N(w_matrix[723]), .A1N(n5156), 
        .Y(n2712) );
  OAI2BB2X1 U6562 ( .B0(n5039), .B1(n5540), .A0N(w_matrix[787]), .A1N(n5165), 
        .Y(n2648) );
  OAI2BB2X1 U6563 ( .B0(n5039), .B1(n5575), .A0N(w_matrix[915]), .A1N(n5173), 
        .Y(n2520) );
  OAI2BB2X1 U6564 ( .B0(n5038), .B1(n5461), .A0N(w_matrix[321]), .A1N(n5120), 
        .Y(n3114) );
  OAI2BB2X1 U6565 ( .B0(n5038), .B1(n5483), .A0N(w_matrix[449]), .A1N(n5136), 
        .Y(n2986) );
  OAI2BB2X1 U6566 ( .B0(n5038), .B1(n5538), .A0N(w_matrix[769]), .A1N(n5164), 
        .Y(n2666) );
  OAI2BB2X1 U6567 ( .B0(n5038), .B1(n5573), .A0N(w_matrix[897]), .A1N(n5172), 
        .Y(n2538) );
  OAI2BB2X1 U6568 ( .B0(n5037), .B1(n5408), .A0N(w_matrix[20]), .A1N(n5093), 
        .Y(n3415) );
  OAI2BB2X1 U6569 ( .B0(n5037), .B1(n5430), .A0N(w_matrix[148]), .A1N(n5103), 
        .Y(n3287) );
  OAI2BB2X1 U6570 ( .B0(n5037), .B1(n5453), .A0N(w_matrix[276]), .A1N(n5113), 
        .Y(n3159) );
  OAI2BB2X1 U6571 ( .B0(n5037), .B1(n5463), .A0N(w_matrix[340]), .A1N(n5121), 
        .Y(n3095) );
  OAI2BB2X1 U6572 ( .B0(n5037), .B1(n5475), .A0N(w_matrix[404]), .A1N(n5129), 
        .Y(n3031) );
  OAI2BB2X1 U6573 ( .B0(n5037), .B1(n5485), .A0N(w_matrix[468]), .A1N(n5137), 
        .Y(n2967) );
  OAI2BB2X1 U6574 ( .B0(n5037), .B1(n5507), .A0N(w_matrix[596]), .A1N(n5145), 
        .Y(n2839) );
  OAI2BB2X1 U6575 ( .B0(n5037), .B1(n5530), .A0N(w_matrix[724]), .A1N(n5156), 
        .Y(n2711) );
  OAI2BB2X1 U6576 ( .B0(n5037), .B1(n5540), .A0N(w_matrix[788]), .A1N(n5165), 
        .Y(n2647) );
  OAI2BB2X1 U6577 ( .B0(n5037), .B1(n5575), .A0N(w_matrix[916]), .A1N(n5173), 
        .Y(n2519) );
  OAI2BB2X1 U6578 ( .B0(n5036), .B1(n5408), .A0N(w_matrix[21]), .A1N(n5093), 
        .Y(n3414) );
  OAI2BB2X1 U6579 ( .B0(n5036), .B1(n5430), .A0N(w_matrix[149]), .A1N(n5103), 
        .Y(n3286) );
  OAI2BB2X1 U6580 ( .B0(n5036), .B1(n5453), .A0N(w_matrix[277]), .A1N(n5113), 
        .Y(n3158) );
  OAI2BB2X1 U6581 ( .B0(n5036), .B1(n5462), .A0N(w_matrix[341]), .A1N(n5121), 
        .Y(n3094) );
  OAI2BB2X1 U6582 ( .B0(n5036), .B1(n5475), .A0N(w_matrix[405]), .A1N(n5129), 
        .Y(n3030) );
  OAI2BB2X1 U6583 ( .B0(n5036), .B1(n5484), .A0N(w_matrix[469]), .A1N(n5137), 
        .Y(n2966) );
  OAI2BB2X1 U6584 ( .B0(n5036), .B1(n5507), .A0N(w_matrix[597]), .A1N(n5145), 
        .Y(n2838) );
  OAI2BB2X1 U6585 ( .B0(n5036), .B1(n5525), .A0N(w_matrix[725]), .A1N(n5156), 
        .Y(n2710) );
  OAI2BB2X1 U6586 ( .B0(n5036), .B1(n5539), .A0N(w_matrix[789]), .A1N(n5165), 
        .Y(n2646) );
  OAI2BB2X1 U6587 ( .B0(n5036), .B1(n5574), .A0N(w_matrix[917]), .A1N(n5173), 
        .Y(n2518) );
  OAI2BB2X1 U6588 ( .B0(n5035), .B1(n5409), .A0N(w_matrix[22]), .A1N(n5094), 
        .Y(n3413) );
  OAI2BB2X1 U6589 ( .B0(n5035), .B1(n5431), .A0N(w_matrix[150]), .A1N(n5104), 
        .Y(n3285) );
  OAI2BB2X1 U6590 ( .B0(n5035), .B1(n5453), .A0N(w_matrix[278]), .A1N(n5113), 
        .Y(n3157) );
  OAI2BB2X1 U6591 ( .B0(n5035), .B1(n5463), .A0N(w_matrix[342]), .A1N(n5121), 
        .Y(n3093) );
  OAI2BB2X1 U6592 ( .B0(n5035), .B1(n5475), .A0N(w_matrix[406]), .A1N(n5129), 
        .Y(n3029) );
  OAI2BB2X1 U6593 ( .B0(n5035), .B1(n5485), .A0N(w_matrix[470]), .A1N(n5137), 
        .Y(n2965) );
  OAI2BB2X1 U6594 ( .B0(n5035), .B1(n5508), .A0N(w_matrix[598]), .A1N(n5146), 
        .Y(n2837) );
  OAI2BB2X1 U6595 ( .B0(n5035), .B1(n5530), .A0N(w_matrix[726]), .A1N(n5157), 
        .Y(n2709) );
  OAI2BB2X1 U6596 ( .B0(n5035), .B1(n5540), .A0N(w_matrix[790]), .A1N(n5165), 
        .Y(n2645) );
  OAI2BB2X1 U6597 ( .B0(n5035), .B1(n5575), .A0N(w_matrix[918]), .A1N(n5173), 
        .Y(n2517) );
  OAI2BB2X1 U6598 ( .B0(n5034), .B1(n5409), .A0N(w_matrix[23]), .A1N(n5094), 
        .Y(n3412) );
  OAI2BB2X1 U6599 ( .B0(n5034), .B1(n5431), .A0N(w_matrix[151]), .A1N(n5104), 
        .Y(n3284) );
  OAI2BB2X1 U6600 ( .B0(n5034), .B1(n5453), .A0N(w_matrix[279]), .A1N(n5113), 
        .Y(n3156) );
  OAI2BB2X1 U6601 ( .B0(n5034), .B1(n5462), .A0N(w_matrix[343]), .A1N(n5121), 
        .Y(n3092) );
  OAI2BB2X1 U6602 ( .B0(n5034), .B1(n5475), .A0N(w_matrix[407]), .A1N(n5129), 
        .Y(n3028) );
  OAI2BB2X1 U6603 ( .B0(n5034), .B1(n5484), .A0N(w_matrix[471]), .A1N(n5137), 
        .Y(n2964) );
  OAI2BB2X1 U6604 ( .B0(n5034), .B1(n5508), .A0N(w_matrix[599]), .A1N(n5146), 
        .Y(n2836) );
  OAI2BB2X1 U6605 ( .B0(n5034), .B1(n5530), .A0N(w_matrix[727]), .A1N(n5157), 
        .Y(n2708) );
  OAI2BB2X1 U6606 ( .B0(n5034), .B1(n5539), .A0N(w_matrix[791]), .A1N(n5165), 
        .Y(n2644) );
  OAI2BB2X1 U6607 ( .B0(n5034), .B1(n5574), .A0N(w_matrix[919]), .A1N(n5173), 
        .Y(n2516) );
  OAI2BB2X1 U6608 ( .B0(n5033), .B1(n5409), .A0N(w_matrix[24]), .A1N(n5094), 
        .Y(n3411) );
  OAI2BB2X1 U6609 ( .B0(n5033), .B1(n5431), .A0N(w_matrix[152]), .A1N(n5104), 
        .Y(n3283) );
  OAI2BB2X1 U6610 ( .B0(n5033), .B1(n5452), .A0N(w_matrix[280]), .A1N(n5113), 
        .Y(n3155) );
  OAI2BB2X1 U6611 ( .B0(n5033), .B1(n5462), .A0N(w_matrix[344]), .A1N(n5121), 
        .Y(n3091) );
  OAI2BB2X1 U6612 ( .B0(n5033), .B1(n5474), .A0N(w_matrix[408]), .A1N(n5129), 
        .Y(n3027) );
  OAI2BB2X1 U6613 ( .B0(n5033), .B1(n5484), .A0N(w_matrix[472]), .A1N(n5137), 
        .Y(n2963) );
  OAI2BB2X1 U6614 ( .B0(n5033), .B1(n5508), .A0N(w_matrix[600]), .A1N(n5146), 
        .Y(n2835) );
  OAI2BB2X1 U6615 ( .B0(n5033), .B1(n5530), .A0N(w_matrix[728]), .A1N(n5157), 
        .Y(n2707) );
  OAI2BB2X1 U6616 ( .B0(n5033), .B1(n5539), .A0N(w_matrix[792]), .A1N(n5165), 
        .Y(n2643) );
  OAI2BB2X1 U6617 ( .B0(n5033), .B1(n5574), .A0N(w_matrix[920]), .A1N(n5173), 
        .Y(n2515) );
  OAI2BB2X1 U6618 ( .B0(n5032), .B1(n5409), .A0N(w_matrix[25]), .A1N(n5094), 
        .Y(n3410) );
  OAI2BB2X1 U6619 ( .B0(n5032), .B1(n5431), .A0N(w_matrix[153]), .A1N(n5104), 
        .Y(n3282) );
  OAI2BB2X1 U6620 ( .B0(n5032), .B1(n5452), .A0N(w_matrix[281]), .A1N(n5113), 
        .Y(n3154) );
  OAI2BB2X1 U6621 ( .B0(n5032), .B1(n5461), .A0N(w_matrix[345]), .A1N(n5121), 
        .Y(n3090) );
  OAI2BB2X1 U6622 ( .B0(n5032), .B1(n5474), .A0N(w_matrix[409]), .A1N(n5129), 
        .Y(n3026) );
  OAI2BB2X1 U6623 ( .B0(n5032), .B1(n5483), .A0N(w_matrix[473]), .A1N(n5137), 
        .Y(n2962) );
  OAI2BB2X1 U6624 ( .B0(n5032), .B1(n5508), .A0N(w_matrix[601]), .A1N(n5146), 
        .Y(n2834) );
  OAI2BB2X1 U6625 ( .B0(n5032), .B1(n5530), .A0N(w_matrix[729]), .A1N(n5157), 
        .Y(n2706) );
  OAI2BB2X1 U6626 ( .B0(n5032), .B1(n5538), .A0N(w_matrix[793]), .A1N(n5165), 
        .Y(n2642) );
  OAI2BB2X1 U6627 ( .B0(n5032), .B1(n5573), .A0N(w_matrix[921]), .A1N(n5173), 
        .Y(n2514) );
  OAI2BB2X1 U6628 ( .B0(n5031), .B1(n5409), .A0N(w_matrix[26]), .A1N(n5094), 
        .Y(n3409) );
  OAI2BB2X1 U6629 ( .B0(n5031), .B1(n5431), .A0N(w_matrix[154]), .A1N(n5104), 
        .Y(n3281) );
  OAI2BB2X1 U6630 ( .B0(n5031), .B1(n5452), .A0N(w_matrix[282]), .A1N(n5114), 
        .Y(n3153) );
  OAI2BB2X1 U6631 ( .B0(n5031), .B1(n5463), .A0N(w_matrix[346]), .A1N(n5122), 
        .Y(n3089) );
  OAI2BB2X1 U6632 ( .B0(n5031), .B1(n5474), .A0N(w_matrix[410]), .A1N(n5130), 
        .Y(n3025) );
  OAI2BB2X1 U6633 ( .B0(n5031), .B1(n5485), .A0N(w_matrix[474]), .A1N(n5138), 
        .Y(n2961) );
  OAI2BB2X1 U6634 ( .B0(n5031), .B1(n5508), .A0N(w_matrix[602]), .A1N(n5146), 
        .Y(n2833) );
  OAI2BB2X1 U6635 ( .B0(n5031), .B1(n5530), .A0N(w_matrix[730]), .A1N(n5157), 
        .Y(n2705) );
  OAI2BB2X1 U6636 ( .B0(n5031), .B1(n5540), .A0N(w_matrix[794]), .A1N(n5166), 
        .Y(n2641) );
  OAI2BB2X1 U6637 ( .B0(n5031), .B1(n5575), .A0N(w_matrix[922]), .A1N(n5174), 
        .Y(n2513) );
  OAI2BB2X1 U6638 ( .B0(n5030), .B1(n5409), .A0N(w_matrix[27]), .A1N(n5094), 
        .Y(n3408) );
  OAI2BB2X1 U6639 ( .B0(n5030), .B1(n5431), .A0N(w_matrix[155]), .A1N(n5104), 
        .Y(n3280) );
  OAI2BB2X1 U6640 ( .B0(n5030), .B1(n5452), .A0N(w_matrix[283]), .A1N(n5114), 
        .Y(n3152) );
  OAI2BB2X1 U6641 ( .B0(n5030), .B1(n5462), .A0N(w_matrix[347]), .A1N(n5122), 
        .Y(n3088) );
  OAI2BB2X1 U6642 ( .B0(n5030), .B1(n5474), .A0N(w_matrix[411]), .A1N(n5130), 
        .Y(n3024) );
  OAI2BB2X1 U6643 ( .B0(n5030), .B1(n5484), .A0N(w_matrix[475]), .A1N(n5138), 
        .Y(n2960) );
  OAI2BB2X1 U6644 ( .B0(n5030), .B1(n5508), .A0N(w_matrix[603]), .A1N(n5146), 
        .Y(n2832) );
  OAI2BB2X1 U6645 ( .B0(n5030), .B1(n5530), .A0N(w_matrix[731]), .A1N(n5157), 
        .Y(n2704) );
  OAI2BB2X1 U6646 ( .B0(n5030), .B1(n5539), .A0N(w_matrix[795]), .A1N(n5166), 
        .Y(n2640) );
  OAI2BB2X1 U6647 ( .B0(n5030), .B1(n5574), .A0N(w_matrix[923]), .A1N(n5174), 
        .Y(n2512) );
  OAI2BB2X1 U6648 ( .B0(n5029), .B1(n5409), .A0N(w_matrix[28]), .A1N(n5094), 
        .Y(n3407) );
  OAI2BB2X1 U6649 ( .B0(n5029), .B1(n5431), .A0N(w_matrix[156]), .A1N(n5104), 
        .Y(n3279) );
  OAI2BB2X1 U6650 ( .B0(n5029), .B1(n5452), .A0N(w_matrix[284]), .A1N(n5114), 
        .Y(n3151) );
  OAI2BB2X1 U6651 ( .B0(n5029), .B1(n5463), .A0N(w_matrix[348]), .A1N(n5122), 
        .Y(n3087) );
  OAI2BB2X1 U6652 ( .B0(n5029), .B1(n5474), .A0N(w_matrix[412]), .A1N(n5130), 
        .Y(n3023) );
  OAI2BB2X1 U6653 ( .B0(n5029), .B1(n5485), .A0N(w_matrix[476]), .A1N(n5138), 
        .Y(n2959) );
  OAI2BB2X1 U6654 ( .B0(n5029), .B1(n5508), .A0N(w_matrix[604]), .A1N(n5146), 
        .Y(n2831) );
  OAI2BB2X1 U6655 ( .B0(n5029), .B1(n5530), .A0N(w_matrix[732]), .A1N(n5157), 
        .Y(n2703) );
  OAI2BB2X1 U6656 ( .B0(n5029), .B1(n5540), .A0N(w_matrix[796]), .A1N(n5166), 
        .Y(n2639) );
  OAI2BB2X1 U6657 ( .B0(n5029), .B1(n5575), .A0N(w_matrix[924]), .A1N(n5174), 
        .Y(n2511) );
  OAI2BB2X1 U6658 ( .B0(n5028), .B1(n5409), .A0N(w_matrix[29]), .A1N(n5094), 
        .Y(n3406) );
  OAI2BB2X1 U6659 ( .B0(n5028), .B1(n5431), .A0N(w_matrix[157]), .A1N(n5104), 
        .Y(n3278) );
  OAI2BB2X1 U6660 ( .B0(n5028), .B1(n5452), .A0N(w_matrix[285]), .A1N(n5114), 
        .Y(n3150) );
  OAI2BB2X1 U6661 ( .B0(n5028), .B1(n5463), .A0N(w_matrix[349]), .A1N(n5122), 
        .Y(n3086) );
  OAI2BB2X1 U6662 ( .B0(n5028), .B1(n5474), .A0N(w_matrix[413]), .A1N(n5130), 
        .Y(n3022) );
  OAI2BB2X1 U6663 ( .B0(n5028), .B1(n5485), .A0N(w_matrix[477]), .A1N(n5138), 
        .Y(n2958) );
  OAI2BB2X1 U6664 ( .B0(n5028), .B1(n5508), .A0N(w_matrix[605]), .A1N(n5146), 
        .Y(n2830) );
  OAI2BB2X1 U6665 ( .B0(n5028), .B1(n5530), .A0N(w_matrix[733]), .A1N(n5157), 
        .Y(n2702) );
  OAI2BB2X1 U6666 ( .B0(n5028), .B1(n5540), .A0N(w_matrix[797]), .A1N(n5166), 
        .Y(n2638) );
  OAI2BB2X1 U6667 ( .B0(n5028), .B1(n5575), .A0N(w_matrix[925]), .A1N(n5174), 
        .Y(n2510) );
  OAI2BB2X1 U6668 ( .B0(n5027), .B1(n5461), .A0N(w_matrix[322]), .A1N(n5120), 
        .Y(n3113) );
  OAI2BB2X1 U6669 ( .B0(n5027), .B1(n5483), .A0N(w_matrix[450]), .A1N(n5136), 
        .Y(n2985) );
  OAI2BB2X1 U6670 ( .B0(n5027), .B1(n5538), .A0N(w_matrix[770]), .A1N(n5164), 
        .Y(n2665) );
  OAI2BB2X1 U6671 ( .B0(n5027), .B1(n5573), .A0N(w_matrix[898]), .A1N(n5172), 
        .Y(n2537) );
  OAI2BB2X1 U6672 ( .B0(n5026), .B1(n5409), .A0N(w_matrix[30]), .A1N(n5094), 
        .Y(n3405) );
  OAI2BB2X1 U6673 ( .B0(n5026), .B1(n5431), .A0N(w_matrix[158]), .A1N(n5104), 
        .Y(n3277) );
  OAI2BB2X1 U6674 ( .B0(n5026), .B1(n5452), .A0N(w_matrix[286]), .A1N(n5114), 
        .Y(n3149) );
  OAI2BB2X1 U6675 ( .B0(n5026), .B1(n5463), .A0N(w_matrix[350]), .A1N(n5122), 
        .Y(n3085) );
  OAI2BB2X1 U6676 ( .B0(n5026), .B1(n5474), .A0N(w_matrix[414]), .A1N(n5130), 
        .Y(n3021) );
  OAI2BB2X1 U6677 ( .B0(n5026), .B1(n5485), .A0N(w_matrix[478]), .A1N(n5138), 
        .Y(n2957) );
  OAI2BB2X1 U6678 ( .B0(n5026), .B1(n5508), .A0N(w_matrix[606]), .A1N(n5146), 
        .Y(n2829) );
  OAI2BB2X1 U6679 ( .B0(n5026), .B1(n5530), .A0N(w_matrix[734]), .A1N(n5157), 
        .Y(n2701) );
  OAI2BB2X1 U6680 ( .B0(n5026), .B1(n5540), .A0N(w_matrix[798]), .A1N(n5166), 
        .Y(n2637) );
  OAI2BB2X1 U6681 ( .B0(n5026), .B1(n5575), .A0N(w_matrix[926]), .A1N(n5174), 
        .Y(n2509) );
  OAI2BB2X1 U6682 ( .B0(n5025), .B1(n5409), .A0N(w_matrix[31]), .A1N(n5094), 
        .Y(n3404) );
  OAI2BB2X1 U6683 ( .B0(n5025), .B1(n5431), .A0N(w_matrix[159]), .A1N(n5104), 
        .Y(n3276) );
  OAI2BB2X1 U6684 ( .B0(n5025), .B1(n5452), .A0N(w_matrix[287]), .A1N(n5114), 
        .Y(n3148) );
  OAI2BB2X1 U6685 ( .B0(n5025), .B1(n5461), .A0N(w_matrix[351]), .A1N(n5122), 
        .Y(n3084) );
  OAI2BB2X1 U6686 ( .B0(n5025), .B1(n5474), .A0N(w_matrix[415]), .A1N(n5130), 
        .Y(n3020) );
  OAI2BB2X1 U6687 ( .B0(n5025), .B1(n5483), .A0N(w_matrix[479]), .A1N(n5138), 
        .Y(n2956) );
  OAI2BB2X1 U6688 ( .B0(n5025), .B1(n5508), .A0N(w_matrix[607]), .A1N(n5146), 
        .Y(n2828) );
  OAI2BB2X1 U6689 ( .B0(n5025), .B1(n5530), .A0N(w_matrix[735]), .A1N(n5157), 
        .Y(n2700) );
  OAI2BB2X1 U6690 ( .B0(n5025), .B1(n5538), .A0N(w_matrix[799]), .A1N(n5166), 
        .Y(n2636) );
  OAI2BB2X1 U6691 ( .B0(n5025), .B1(n5573), .A0N(w_matrix[927]), .A1N(n5174), 
        .Y(n2508) );
  OAI2BB2X1 U6692 ( .B0(n5024), .B1(n5409), .A0N(w_matrix[32]), .A1N(n5094), 
        .Y(n3403) );
  OAI2BB2X1 U6693 ( .B0(n5024), .B1(n5431), .A0N(w_matrix[160]), .A1N(n5104), 
        .Y(n3275) );
  OAI2BB2X1 U6694 ( .B0(n5024), .B1(n5452), .A0N(w_matrix[288]), .A1N(n5114), 
        .Y(n3147) );
  OAI2BB2X1 U6695 ( .B0(n5024), .B1(n5464), .A0N(w_matrix[352]), .A1N(n5122), 
        .Y(n3083) );
  OAI2BB2X1 U6696 ( .B0(n5024), .B1(n5474), .A0N(w_matrix[416]), .A1N(n5130), 
        .Y(n3019) );
  OAI2BB2X1 U6697 ( .B0(n5024), .B1(n5486), .A0N(w_matrix[480]), .A1N(n5138), 
        .Y(n2955) );
  OAI2BB2X1 U6698 ( .B0(n5024), .B1(n5508), .A0N(w_matrix[608]), .A1N(n5146), 
        .Y(n2827) );
  OAI2BB2X1 U6699 ( .B0(n5024), .B1(n5530), .A0N(w_matrix[736]), .A1N(n5157), 
        .Y(n2699) );
  OAI2BB2X1 U6700 ( .B0(n5024), .B1(n5541), .A0N(w_matrix[800]), .A1N(n5166), 
        .Y(n2635) );
  OAI2BB2X1 U6701 ( .B0(n5024), .B1(n5576), .A0N(w_matrix[928]), .A1N(n5174), 
        .Y(n2507) );
  OAI2BB2X1 U6702 ( .B0(n5023), .B1(n5409), .A0N(w_matrix[33]), .A1N(n5094), 
        .Y(n3402) );
  OAI2BB2X1 U6703 ( .B0(n5023), .B1(n5431), .A0N(w_matrix[161]), .A1N(n5104), 
        .Y(n3274) );
  OAI2BB2X1 U6704 ( .B0(n5023), .B1(n5452), .A0N(w_matrix[289]), .A1N(n5114), 
        .Y(n3146) );
  OAI2BB2X1 U6705 ( .B0(n5023), .B1(n5463), .A0N(w_matrix[353]), .A1N(n5122), 
        .Y(n3082) );
  OAI2BB2X1 U6706 ( .B0(n5023), .B1(n5474), .A0N(w_matrix[417]), .A1N(n5130), 
        .Y(n3018) );
  OAI2BB2X1 U6707 ( .B0(n5023), .B1(n5485), .A0N(w_matrix[481]), .A1N(n5138), 
        .Y(n2954) );
  OAI2BB2X1 U6708 ( .B0(n5023), .B1(n5508), .A0N(w_matrix[609]), .A1N(n5146), 
        .Y(n2826) );
  OAI2BB2X1 U6709 ( .B0(n5023), .B1(n5530), .A0N(w_matrix[737]), .A1N(n5157), 
        .Y(n2698) );
  OAI2BB2X1 U6710 ( .B0(n5023), .B1(n5540), .A0N(w_matrix[801]), .A1N(n5166), 
        .Y(n2634) );
  OAI2BB2X1 U6711 ( .B0(n5023), .B1(n5575), .A0N(w_matrix[929]), .A1N(n5174), 
        .Y(n2506) );
  OAI2BB2X1 U6712 ( .B0(n5022), .B1(n5409), .A0N(w_matrix[34]), .A1N(n5094), 
        .Y(n3401) );
  OAI2BB2X1 U6713 ( .B0(n5022), .B1(n5431), .A0N(w_matrix[162]), .A1N(n5104), 
        .Y(n3273) );
  OAI2BB2X1 U6714 ( .B0(n5022), .B1(n5452), .A0N(w_matrix[290]), .A1N(n5114), 
        .Y(n3145) );
  OAI2BB2X1 U6715 ( .B0(n5022), .B1(n5464), .A0N(w_matrix[354]), .A1N(n5122), 
        .Y(n3081) );
  OAI2BB2X1 U6716 ( .B0(n5022), .B1(n5474), .A0N(w_matrix[418]), .A1N(n5130), 
        .Y(n3017) );
  OAI2BB2X1 U6717 ( .B0(n5022), .B1(n5486), .A0N(w_matrix[482]), .A1N(n5138), 
        .Y(n2953) );
  OAI2BB2X1 U6718 ( .B0(n5022), .B1(n5508), .A0N(w_matrix[610]), .A1N(n5146), 
        .Y(n2825) );
  OAI2BB2X1 U6719 ( .B0(n5022), .B1(n5530), .A0N(w_matrix[738]), .A1N(n5157), 
        .Y(n2697) );
  OAI2BB2X1 U6720 ( .B0(n5022), .B1(n5541), .A0N(w_matrix[802]), .A1N(n5166), 
        .Y(n2633) );
  OAI2BB2X1 U6721 ( .B0(n5022), .B1(n5576), .A0N(w_matrix[930]), .A1N(n5174), 
        .Y(n2505) );
  OAI2BB2X1 U6722 ( .B0(n5021), .B1(n5410), .A0N(w_matrix[35]), .A1N(n5095), 
        .Y(n3400) );
  OAI2BB2X1 U6723 ( .B0(n5021), .B1(n5432), .A0N(w_matrix[163]), .A1N(n5105), 
        .Y(n3272) );
  OAI2BB2X1 U6724 ( .B0(n5021), .B1(n5452), .A0N(w_matrix[291]), .A1N(n5114), 
        .Y(n3144) );
  OAI2BB2X1 U6725 ( .B0(n5021), .B1(n5464), .A0N(w_matrix[355]), .A1N(n5122), 
        .Y(n3080) );
  OAI2BB2X1 U6726 ( .B0(n5021), .B1(n5474), .A0N(w_matrix[419]), .A1N(n5130), 
        .Y(n3016) );
  OAI2BB2X1 U6727 ( .B0(n5021), .B1(n5486), .A0N(w_matrix[483]), .A1N(n5138), 
        .Y(n2952) );
  OAI2BB2X1 U6728 ( .B0(n5021), .B1(n5509), .A0N(w_matrix[611]), .A1N(n5147), 
        .Y(n2824) );
  OAI2BB2X1 U6729 ( .B0(n5021), .B1(n5531), .A0N(w_matrix[739]), .A1N(n5158), 
        .Y(n2696) );
  OAI2BB2X1 U6730 ( .B0(n5021), .B1(n5541), .A0N(w_matrix[803]), .A1N(n5166), 
        .Y(n2632) );
  OAI2BB2X1 U6731 ( .B0(n5021), .B1(n5576), .A0N(w_matrix[931]), .A1N(n5174), 
        .Y(n2504) );
  OAI2BB2X1 U6732 ( .B0(n5020), .B1(n5410), .A0N(w_matrix[36]), .A1N(n5095), 
        .Y(n3399) );
  OAI2BB2X1 U6733 ( .B0(n5020), .B1(n5432), .A0N(w_matrix[164]), .A1N(n5105), 
        .Y(n3271) );
  OAI2BB2X1 U6734 ( .B0(n5020), .B1(n5452), .A0N(w_matrix[292]), .A1N(n5114), 
        .Y(n3143) );
  OAI2BB2X1 U6735 ( .B0(n5020), .B1(n5463), .A0N(w_matrix[356]), .A1N(n5122), 
        .Y(n3079) );
  OAI2BB2X1 U6736 ( .B0(n5020), .B1(n5474), .A0N(w_matrix[420]), .A1N(n5130), 
        .Y(n3015) );
  OAI2BB2X1 U6737 ( .B0(n5020), .B1(n5485), .A0N(w_matrix[484]), .A1N(n5138), 
        .Y(n2951) );
  OAI2BB2X1 U6738 ( .B0(n5020), .B1(n5509), .A0N(w_matrix[612]), .A1N(n5147), 
        .Y(n2823) );
  OAI2BB2X1 U6739 ( .B0(n5020), .B1(n5531), .A0N(w_matrix[740]), .A1N(n5158), 
        .Y(n2695) );
  OAI2BB2X1 U6740 ( .B0(n5020), .B1(n5540), .A0N(w_matrix[804]), .A1N(n5166), 
        .Y(n2631) );
  OAI2BB2X1 U6741 ( .B0(n5020), .B1(n5575), .A0N(w_matrix[932]), .A1N(n5174), 
        .Y(n2503) );
  OAI2BB2X1 U6742 ( .B0(n5019), .B1(n5410), .A0N(w_matrix[37]), .A1N(n5095), 
        .Y(n3398) );
  OAI2BB2X1 U6743 ( .B0(n5019), .B1(n5432), .A0N(w_matrix[165]), .A1N(n5105), 
        .Y(n3270) );
  OAI2BB2X1 U6744 ( .B0(n5019), .B1(n5451), .A0N(w_matrix[293]), .A1N(n5114), 
        .Y(n3142) );
  OAI2BB2X1 U6745 ( .B0(n5019), .B1(n5464), .A0N(w_matrix[357]), .A1N(n5122), 
        .Y(n3078) );
  OAI2BB2X1 U6746 ( .B0(n5019), .B1(n5473), .A0N(w_matrix[421]), .A1N(n5130), 
        .Y(n3014) );
  OAI2BB2X1 U6747 ( .B0(n5019), .B1(n5486), .A0N(w_matrix[485]), .A1N(n5138), 
        .Y(n2950) );
  OAI2BB2X1 U6748 ( .B0(n5019), .B1(n5509), .A0N(w_matrix[613]), .A1N(n5147), 
        .Y(n2822) );
  OAI2BB2X1 U6749 ( .B0(n5019), .B1(n5531), .A0N(w_matrix[741]), .A1N(n5158), 
        .Y(n2694) );
  OAI2BB2X1 U6750 ( .B0(n5019), .B1(n5541), .A0N(w_matrix[805]), .A1N(n5166), 
        .Y(n2630) );
  OAI2BB2X1 U6751 ( .B0(n5019), .B1(n5576), .A0N(w_matrix[933]), .A1N(n5174), 
        .Y(n2502) );
  OAI2BB2X1 U6752 ( .B0(n5018), .B1(n5410), .A0N(w_matrix[38]), .A1N(n5095), 
        .Y(n3397) );
  OAI2BB2X1 U6753 ( .B0(n5018), .B1(n5432), .A0N(w_matrix[166]), .A1N(n5105), 
        .Y(n3269) );
  OAI2BB2X1 U6754 ( .B0(n5018), .B1(n5451), .A0N(w_matrix[294]), .A1N(n5114), 
        .Y(n3141) );
  OAI2BB2X1 U6755 ( .B0(n5018), .B1(n5464), .A0N(w_matrix[358]), .A1N(n5122), 
        .Y(n3077) );
  OAI2BB2X1 U6756 ( .B0(n5018), .B1(n5473), .A0N(w_matrix[422]), .A1N(n5130), 
        .Y(n3013) );
  OAI2BB2X1 U6757 ( .B0(n5018), .B1(n5486), .A0N(w_matrix[486]), .A1N(n5138), 
        .Y(n2949) );
  OAI2BB2X1 U6758 ( .B0(n5018), .B1(n5509), .A0N(w_matrix[614]), .A1N(n5147), 
        .Y(n2821) );
  OAI2BB2X1 U6759 ( .B0(n5018), .B1(n5531), .A0N(w_matrix[742]), .A1N(n5158), 
        .Y(n2693) );
  OAI2BB2X1 U6760 ( .B0(n5018), .B1(n5541), .A0N(w_matrix[806]), .A1N(n5166), 
        .Y(n2629) );
  OAI2BB2X1 U6761 ( .B0(n5018), .B1(n5576), .A0N(w_matrix[934]), .A1N(n5174), 
        .Y(n2501) );
  OAI2BB2X1 U6762 ( .B0(n5017), .B1(n5410), .A0N(w_matrix[39]), .A1N(n5095), 
        .Y(n3396) );
  OAI2BB2X1 U6763 ( .B0(n5017), .B1(n5432), .A0N(w_matrix[167]), .A1N(n5105), 
        .Y(n3268) );
  OAI2BB2X1 U6764 ( .B0(n5017), .B1(n5451), .A0N(w_matrix[295]), .A1N(n5115), 
        .Y(n3140) );
  OAI2BB2X1 U6765 ( .B0(n5017), .B1(n5463), .A0N(w_matrix[359]), .A1N(n5123), 
        .Y(n3076) );
  OAI2BB2X1 U6766 ( .B0(n5017), .B1(n5473), .A0N(w_matrix[423]), .A1N(n5131), 
        .Y(n3012) );
  OAI2BB2X1 U6767 ( .B0(n5017), .B1(n5485), .A0N(w_matrix[487]), .A1N(n5139), 
        .Y(n2948) );
  OAI2BB2X1 U6768 ( .B0(n5017), .B1(n5509), .A0N(w_matrix[615]), .A1N(n5147), 
        .Y(n2820) );
  OAI2BB2X1 U6769 ( .B0(n5017), .B1(n5531), .A0N(w_matrix[743]), .A1N(n5158), 
        .Y(n2692) );
  OAI2BB2X1 U6770 ( .B0(n5017), .B1(n5540), .A0N(w_matrix[807]), .A1N(n5167), 
        .Y(n2628) );
  OAI2BB2X1 U6771 ( .B0(n5017), .B1(n5575), .A0N(w_matrix[935]), .A1N(n5175), 
        .Y(n2500) );
  OAI2BB2X1 U6772 ( .B0(n5016), .B1(n5461), .A0N(w_matrix[323]), .A1N(n5120), 
        .Y(n3112) );
  OAI2BB2X1 U6773 ( .B0(n5016), .B1(n5483), .A0N(w_matrix[451]), .A1N(n5136), 
        .Y(n2984) );
  OAI2BB2X1 U6774 ( .B0(n5016), .B1(n5538), .A0N(w_matrix[771]), .A1N(n5164), 
        .Y(n2664) );
  OAI2BB2X1 U6775 ( .B0(n5016), .B1(n5573), .A0N(w_matrix[899]), .A1N(n5172), 
        .Y(n2536) );
  OAI2BB2X1 U6776 ( .B0(n5015), .B1(n5410), .A0N(w_matrix[40]), .A1N(n5095), 
        .Y(n3395) );
  OAI2BB2X1 U6777 ( .B0(n5015), .B1(n5432), .A0N(w_matrix[168]), .A1N(n5105), 
        .Y(n3267) );
  OAI2BB2X1 U6778 ( .B0(n5015), .B1(n5451), .A0N(w_matrix[296]), .A1N(n5115), 
        .Y(n3139) );
  OAI2BB2X1 U6779 ( .B0(n5015), .B1(n5464), .A0N(w_matrix[360]), .A1N(n5123), 
        .Y(n3075) );
  OAI2BB2X1 U6780 ( .B0(n5015), .B1(n5473), .A0N(w_matrix[424]), .A1N(n5131), 
        .Y(n3011) );
  OAI2BB2X1 U6781 ( .B0(n5015), .B1(n5486), .A0N(w_matrix[488]), .A1N(n5139), 
        .Y(n2947) );
  OAI2BB2X1 U6782 ( .B0(n5015), .B1(n5509), .A0N(w_matrix[616]), .A1N(n5147), 
        .Y(n2819) );
  OAI2BB2X1 U6783 ( .B0(n5015), .B1(n5531), .A0N(w_matrix[744]), .A1N(n5158), 
        .Y(n2691) );
  OAI2BB2X1 U6784 ( .B0(n5015), .B1(n5541), .A0N(w_matrix[808]), .A1N(n5167), 
        .Y(n2627) );
  OAI2BB2X1 U6785 ( .B0(n5015), .B1(n5576), .A0N(w_matrix[936]), .A1N(n5175), 
        .Y(n2499) );
  OAI2BB2X1 U6786 ( .B0(n5014), .B1(n5410), .A0N(w_matrix[41]), .A1N(n5095), 
        .Y(n3394) );
  OAI2BB2X1 U6787 ( .B0(n5014), .B1(n5432), .A0N(w_matrix[169]), .A1N(n5105), 
        .Y(n3266) );
  OAI2BB2X1 U6788 ( .B0(n5014), .B1(n5451), .A0N(w_matrix[297]), .A1N(n5115), 
        .Y(n3138) );
  OAI2BB2X1 U6789 ( .B0(n5014), .B1(n5464), .A0N(w_matrix[361]), .A1N(n5123), 
        .Y(n3074) );
  OAI2BB2X1 U6790 ( .B0(n5014), .B1(n5473), .A0N(w_matrix[425]), .A1N(n5131), 
        .Y(n3010) );
  OAI2BB2X1 U6791 ( .B0(n5014), .B1(n5486), .A0N(w_matrix[489]), .A1N(n5139), 
        .Y(n2946) );
  OAI2BB2X1 U6792 ( .B0(n5014), .B1(n5509), .A0N(w_matrix[617]), .A1N(n5147), 
        .Y(n2818) );
  OAI2BB2X1 U6793 ( .B0(n5014), .B1(n5531), .A0N(w_matrix[745]), .A1N(n5158), 
        .Y(n2690) );
  OAI2BB2X1 U6794 ( .B0(n5014), .B1(n5541), .A0N(w_matrix[809]), .A1N(n5167), 
        .Y(n2626) );
  OAI2BB2X1 U6795 ( .B0(n5014), .B1(n5576), .A0N(w_matrix[937]), .A1N(n5175), 
        .Y(n2498) );
  OAI2BB2X1 U6796 ( .B0(n5013), .B1(n5410), .A0N(w_matrix[42]), .A1N(n5095), 
        .Y(n3393) );
  OAI2BB2X1 U6797 ( .B0(n5013), .B1(n5432), .A0N(w_matrix[170]), .A1N(n5105), 
        .Y(n3265) );
  OAI2BB2X1 U6798 ( .B0(n5013), .B1(n5451), .A0N(w_matrix[298]), .A1N(n5115), 
        .Y(n3137) );
  OAI2BB2X1 U6799 ( .B0(n5013), .B1(n5463), .A0N(w_matrix[362]), .A1N(n5123), 
        .Y(n3073) );
  OAI2BB2X1 U6800 ( .B0(n5013), .B1(n5473), .A0N(w_matrix[426]), .A1N(n5131), 
        .Y(n3009) );
  OAI2BB2X1 U6801 ( .B0(n5013), .B1(n5485), .A0N(w_matrix[490]), .A1N(n5139), 
        .Y(n2945) );
  OAI2BB2X1 U6802 ( .B0(n5013), .B1(n5509), .A0N(w_matrix[618]), .A1N(n5147), 
        .Y(n2817) );
  OAI2BB2X1 U6803 ( .B0(n5013), .B1(n5531), .A0N(w_matrix[746]), .A1N(n5158), 
        .Y(n2689) );
  OAI2BB2X1 U6804 ( .B0(n5013), .B1(n5540), .A0N(w_matrix[810]), .A1N(n5167), 
        .Y(n2625) );
  OAI2BB2X1 U6805 ( .B0(n5013), .B1(n5575), .A0N(w_matrix[938]), .A1N(n5175), 
        .Y(n2497) );
  OAI2BB2X1 U6806 ( .B0(n5012), .B1(n5410), .A0N(w_matrix[43]), .A1N(n5095), 
        .Y(n3392) );
  OAI2BB2X1 U6807 ( .B0(n5012), .B1(n5432), .A0N(w_matrix[171]), .A1N(n5105), 
        .Y(n3264) );
  OAI2BB2X1 U6808 ( .B0(n5012), .B1(n5451), .A0N(w_matrix[299]), .A1N(n5115), 
        .Y(n3136) );
  OAI2BB2X1 U6809 ( .B0(n5012), .B1(n5464), .A0N(w_matrix[363]), .A1N(n5123), 
        .Y(n3072) );
  OAI2BB2X1 U6810 ( .B0(n5012), .B1(n5473), .A0N(w_matrix[427]), .A1N(n5131), 
        .Y(n3008) );
  OAI2BB2X1 U6811 ( .B0(n5012), .B1(n5486), .A0N(w_matrix[491]), .A1N(n5139), 
        .Y(n2944) );
  OAI2BB2X1 U6812 ( .B0(n5012), .B1(n5509), .A0N(w_matrix[619]), .A1N(n5147), 
        .Y(n2816) );
  OAI2BB2X1 U6813 ( .B0(n5012), .B1(n5531), .A0N(w_matrix[747]), .A1N(n5158), 
        .Y(n2688) );
  OAI2BB2X1 U6814 ( .B0(n5012), .B1(n5541), .A0N(w_matrix[811]), .A1N(n5167), 
        .Y(n2624) );
  OAI2BB2X1 U6815 ( .B0(n5012), .B1(n5576), .A0N(w_matrix[939]), .A1N(n5175), 
        .Y(n2496) );
  OAI2BB2X1 U6816 ( .B0(n5011), .B1(n5410), .A0N(w_matrix[44]), .A1N(n5095), 
        .Y(n3391) );
  OAI2BB2X1 U6817 ( .B0(n5011), .B1(n5432), .A0N(w_matrix[172]), .A1N(n5105), 
        .Y(n3263) );
  OAI2BB2X1 U6818 ( .B0(n5011), .B1(n5451), .A0N(w_matrix[300]), .A1N(n5115), 
        .Y(n3135) );
  OAI2BB2X1 U6819 ( .B0(n5011), .B1(n5463), .A0N(w_matrix[364]), .A1N(n5123), 
        .Y(n3071) );
  OAI2BB2X1 U6820 ( .B0(n5011), .B1(n5473), .A0N(w_matrix[428]), .A1N(n5131), 
        .Y(n3007) );
  OAI2BB2X1 U6821 ( .B0(n5011), .B1(n5485), .A0N(w_matrix[492]), .A1N(n5139), 
        .Y(n2943) );
  OAI2BB2X1 U6822 ( .B0(n5011), .B1(n5509), .A0N(w_matrix[620]), .A1N(n5147), 
        .Y(n2815) );
  OAI2BB2X1 U6823 ( .B0(n5011), .B1(n5531), .A0N(w_matrix[748]), .A1N(n5158), 
        .Y(n2687) );
  OAI2BB2X1 U6824 ( .B0(n5011), .B1(n5540), .A0N(w_matrix[812]), .A1N(n5167), 
        .Y(n2623) );
  OAI2BB2X1 U6825 ( .B0(n5011), .B1(n5575), .A0N(w_matrix[940]), .A1N(n5175), 
        .Y(n2495) );
  OAI2BB2X1 U6826 ( .B0(n5010), .B1(n5410), .A0N(w_matrix[45]), .A1N(n5095), 
        .Y(n3390) );
  OAI2BB2X1 U6827 ( .B0(n5010), .B1(n5432), .A0N(w_matrix[173]), .A1N(n5105), 
        .Y(n3262) );
  OAI2BB2X1 U6828 ( .B0(n5010), .B1(n5451), .A0N(w_matrix[301]), .A1N(n5115), 
        .Y(n3134) );
  OAI2BB2X1 U6829 ( .B0(n5010), .B1(n5464), .A0N(w_matrix[365]), .A1N(n5123), 
        .Y(n3070) );
  OAI2BB2X1 U6830 ( .B0(n5010), .B1(n5473), .A0N(w_matrix[429]), .A1N(n5131), 
        .Y(n3006) );
  OAI2BB2X1 U6831 ( .B0(n5010), .B1(n5486), .A0N(w_matrix[493]), .A1N(n5139), 
        .Y(n2942) );
  OAI2BB2X1 U6832 ( .B0(n5010), .B1(n5509), .A0N(w_matrix[621]), .A1N(n5147), 
        .Y(n2814) );
  OAI2BB2X1 U6833 ( .B0(n5010), .B1(n5531), .A0N(w_matrix[749]), .A1N(n5158), 
        .Y(n2686) );
  OAI2BB2X1 U6834 ( .B0(n5010), .B1(n5541), .A0N(w_matrix[813]), .A1N(n5167), 
        .Y(n2622) );
  OAI2BB2X1 U6835 ( .B0(n5010), .B1(n5576), .A0N(w_matrix[941]), .A1N(n5175), 
        .Y(n2494) );
  OAI2BB2X1 U6836 ( .B0(n5009), .B1(n5410), .A0N(w_matrix[46]), .A1N(n5095), 
        .Y(n3389) );
  OAI2BB2X1 U6837 ( .B0(n5009), .B1(n5432), .A0N(w_matrix[174]), .A1N(n5105), 
        .Y(n3261) );
  OAI2BB2X1 U6838 ( .B0(n5009), .B1(n5451), .A0N(w_matrix[302]), .A1N(n5115), 
        .Y(n3133) );
  OAI2BB2X1 U6839 ( .B0(n5009), .B1(n5473), .A0N(w_matrix[430]), .A1N(n5131), 
        .Y(n3005) );
  OAI2BB2X1 U6840 ( .B0(n5009), .B1(n5509), .A0N(w_matrix[622]), .A1N(n5147), 
        .Y(n2813) );
  OAI2BB2X1 U6841 ( .B0(n5009), .B1(n5531), .A0N(w_matrix[750]), .A1N(n5158), 
        .Y(n2685) );
  OAI2BB2X1 U6842 ( .B0(n5008), .B1(n5410), .A0N(w_matrix[47]), .A1N(n5095), 
        .Y(n3388) );
  OAI2BB2X1 U6843 ( .B0(n5008), .B1(n5432), .A0N(w_matrix[175]), .A1N(n5105), 
        .Y(n3260) );
  OAI2BB2X1 U6844 ( .B0(n5008), .B1(n5451), .A0N(w_matrix[303]), .A1N(n5115), 
        .Y(n3132) );
  OAI2BB2X1 U6845 ( .B0(n5008), .B1(n5464), .A0N(w_matrix[367]), .A1N(n5123), 
        .Y(n3068) );
  OAI2BB2X1 U6846 ( .B0(n5008), .B1(n5473), .A0N(w_matrix[431]), .A1N(n5131), 
        .Y(n3004) );
  OAI2BB2X1 U6847 ( .B0(n5008), .B1(n5486), .A0N(w_matrix[495]), .A1N(n5139), 
        .Y(n2940) );
  OAI2BB2X1 U6848 ( .B0(n5008), .B1(n5509), .A0N(w_matrix[623]), .A1N(n5147), 
        .Y(n2812) );
  OAI2BB2X1 U6849 ( .B0(n5008), .B1(n5531), .A0N(w_matrix[751]), .A1N(n5158), 
        .Y(n2684) );
  OAI2BB2X1 U6850 ( .B0(n5008), .B1(n5541), .A0N(w_matrix[815]), .A1N(n5167), 
        .Y(n2620) );
  OAI2BB2X1 U6851 ( .B0(n5008), .B1(n5576), .A0N(w_matrix[943]), .A1N(n5175), 
        .Y(n2492) );
  OAI2BB2X1 U6852 ( .B0(n5007), .B1(n5411), .A0N(w_matrix[48]), .A1N(n5096), 
        .Y(n3387) );
  OAI2BB2X1 U6853 ( .B0(n5007), .B1(n5433), .A0N(w_matrix[176]), .A1N(n5106), 
        .Y(n3259) );
  OAI2BB2X1 U6854 ( .B0(n5007), .B1(n5451), .A0N(w_matrix[304]), .A1N(n5115), 
        .Y(n3131) );
  OAI2BB2X1 U6855 ( .B0(n5007), .B1(n5464), .A0N(w_matrix[368]), .A1N(n5123), 
        .Y(n3067) );
  OAI2BB2X1 U6856 ( .B0(n5007), .B1(n5473), .A0N(w_matrix[432]), .A1N(n5131), 
        .Y(n3003) );
  OAI2BB2X1 U6857 ( .B0(n5007), .B1(n5486), .A0N(w_matrix[496]), .A1N(n5139), 
        .Y(n2939) );
  OAI2BB2X1 U6858 ( .B0(n5007), .B1(n5510), .A0N(w_matrix[624]), .A1N(n5148), 
        .Y(n2811) );
  OAI2BB2X1 U6859 ( .B0(n5007), .B1(n5532), .A0N(w_matrix[752]), .A1N(n5159), 
        .Y(n2683) );
  OAI2BB2X1 U6860 ( .B0(n5007), .B1(n5541), .A0N(w_matrix[816]), .A1N(n5167), 
        .Y(n2619) );
  OAI2BB2X1 U6861 ( .B0(n5007), .B1(n5576), .A0N(w_matrix[944]), .A1N(n5175), 
        .Y(n2491) );
  OAI2BB2X1 U6862 ( .B0(n5006), .B1(n5411), .A0N(w_matrix[49]), .A1N(n5096), 
        .Y(n3386) );
  OAI2BB2X1 U6863 ( .B0(n5006), .B1(n5433), .A0N(w_matrix[177]), .A1N(n5106), 
        .Y(n3258) );
  OAI2BB2X1 U6864 ( .B0(n5006), .B1(n5451), .A0N(w_matrix[305]), .A1N(n5115), 
        .Y(n3130) );
  OAI2BB2X1 U6865 ( .B0(n5006), .B1(n5473), .A0N(w_matrix[433]), .A1N(n5131), 
        .Y(n3002) );
  OAI2BB2X1 U6866 ( .B0(n5006), .B1(n5510), .A0N(w_matrix[625]), .A1N(n5148), 
        .Y(n2810) );
  OAI2BB2X1 U6867 ( .B0(n5006), .B1(n5532), .A0N(w_matrix[753]), .A1N(n5159), 
        .Y(n2682) );
  OAI2BB2X1 U6868 ( .B0(n5005), .B1(n5461), .A0N(w_matrix[324]), .A1N(n5120), 
        .Y(n3111) );
  OAI2BB2X1 U6869 ( .B0(n5005), .B1(n5483), .A0N(w_matrix[452]), .A1N(n5136), 
        .Y(n2983) );
  OAI2BB2X1 U6870 ( .B0(n5005), .B1(n5538), .A0N(w_matrix[772]), .A1N(n5164), 
        .Y(n2663) );
  OAI2BB2X1 U6871 ( .B0(n5005), .B1(n5573), .A0N(w_matrix[900]), .A1N(n5172), 
        .Y(n2535) );
  OAI2BB2X1 U6872 ( .B0(n5004), .B1(n5411), .A0N(w_matrix[50]), .A1N(n5096), 
        .Y(n3385) );
  OAI2BB2X1 U6873 ( .B0(n5004), .B1(n5433), .A0N(w_matrix[178]), .A1N(n5106), 
        .Y(n3257) );
  OAI2BB2X1 U6874 ( .B0(n5004), .B1(n5450), .A0N(w_matrix[306]), .A1N(n5115), 
        .Y(n3129) );
  OAI2BB2X1 U6875 ( .B0(n5004), .B1(n5472), .A0N(w_matrix[434]), .A1N(n5131), 
        .Y(n3001) );
  OAI2BB2X1 U6876 ( .B0(n5004), .B1(n5510), .A0N(w_matrix[626]), .A1N(n5148), 
        .Y(n2809) );
  OAI2BB2X1 U6877 ( .B0(n5004), .B1(n5532), .A0N(w_matrix[754]), .A1N(n5159), 
        .Y(n2681) );
  OAI2BB2X1 U6878 ( .B0(n5003), .B1(n5411), .A0N(w_matrix[51]), .A1N(n5096), 
        .Y(n3384) );
  OAI2BB2X1 U6879 ( .B0(n5003), .B1(n5433), .A0N(w_matrix[179]), .A1N(n5106), 
        .Y(n3256) );
  OAI2BB2X1 U6880 ( .B0(n5003), .B1(n5450), .A0N(w_matrix[307]), .A1N(n5115), 
        .Y(n3128) );
  OAI2BB2X1 U6881 ( .B0(n5003), .B1(n5464), .A0N(w_matrix[371]), .A1N(n5123), 
        .Y(n3064) );
  OAI2BB2X1 U6882 ( .B0(n5003), .B1(n5472), .A0N(w_matrix[435]), .A1N(n5131), 
        .Y(n3000) );
  OAI2BB2X1 U6883 ( .B0(n5003), .B1(n5486), .A0N(w_matrix[499]), .A1N(n5139), 
        .Y(n2936) );
  OAI2BB2X1 U6884 ( .B0(n5003), .B1(n5510), .A0N(w_matrix[627]), .A1N(n5148), 
        .Y(n2808) );
  OAI2BB2X1 U6885 ( .B0(n5003), .B1(n5532), .A0N(w_matrix[755]), .A1N(n5159), 
        .Y(n2680) );
  OAI2BB2X1 U6886 ( .B0(n5003), .B1(n5541), .A0N(w_matrix[819]), .A1N(n5167), 
        .Y(n2616) );
  OAI2BB2X1 U6887 ( .B0(n5003), .B1(n5576), .A0N(w_matrix[947]), .A1N(n5175), 
        .Y(n2488) );
  OAI2BB2X1 U6888 ( .B0(n5002), .B1(n5411), .A0N(w_matrix[52]), .A1N(n5096), 
        .Y(n3383) );
  OAI2BB2X1 U6889 ( .B0(n5002), .B1(n5433), .A0N(w_matrix[180]), .A1N(n5106), 
        .Y(n3255) );
  OAI2BB2X1 U6890 ( .B0(n5002), .B1(n5450), .A0N(w_matrix[308]), .A1N(n5116), 
        .Y(n3127) );
  OAI2BB2X1 U6891 ( .B0(n5002), .B1(n5472), .A0N(w_matrix[436]), .A1N(n5132), 
        .Y(n2999) );
  OAI2BB2X1 U6892 ( .B0(n5002), .B1(n5510), .A0N(w_matrix[628]), .A1N(n5148), 
        .Y(n2807) );
  OAI2BB2X1 U6893 ( .B0(n5002), .B1(n5532), .A0N(w_matrix[756]), .A1N(n5159), 
        .Y(n2679) );
  OAI2BB2X1 U6894 ( .B0(n5001), .B1(n5411), .A0N(w_matrix[53]), .A1N(n5096), 
        .Y(n3382) );
  OAI2BB2X1 U6895 ( .B0(n5001), .B1(n5433), .A0N(w_matrix[181]), .A1N(n5106), 
        .Y(n3254) );
  OAI2BB2X1 U6896 ( .B0(n5001), .B1(n5450), .A0N(w_matrix[309]), .A1N(n5116), 
        .Y(n3126) );
  OAI2BB2X1 U6897 ( .B0(n5001), .B1(n5472), .A0N(w_matrix[437]), .A1N(n5132), 
        .Y(n2998) );
  OAI2BB2X1 U6898 ( .B0(n5001), .B1(n5510), .A0N(w_matrix[629]), .A1N(n5148), 
        .Y(n2806) );
  OAI2BB2X1 U6899 ( .B0(n5001), .B1(n5532), .A0N(w_matrix[757]), .A1N(n5159), 
        .Y(n2678) );
  OAI2BB2X1 U6900 ( .B0(n5000), .B1(n5411), .A0N(w_matrix[54]), .A1N(n5096), 
        .Y(n3381) );
  OAI2BB2X1 U6901 ( .B0(n5000), .B1(n5433), .A0N(w_matrix[182]), .A1N(n5106), 
        .Y(n3253) );
  OAI2BB2X1 U6902 ( .B0(n5000), .B1(n5450), .A0N(w_matrix[310]), .A1N(n5116), 
        .Y(n3125) );
  OAI2BB2X1 U6903 ( .B0(n5000), .B1(n5464), .A0N(w_matrix[374]), .A1N(n5124), 
        .Y(n3061) );
  OAI2BB2X1 U6904 ( .B0(n5000), .B1(n5472), .A0N(w_matrix[438]), .A1N(n5132), 
        .Y(n2997) );
  OAI2BB2X1 U6905 ( .B0(n5000), .B1(n5486), .A0N(w_matrix[502]), .A1N(n5140), 
        .Y(n2933) );
  OAI2BB2X1 U6906 ( .B0(n5000), .B1(n5510), .A0N(w_matrix[630]), .A1N(n5148), 
        .Y(n2805) );
  OAI2BB2X1 U6907 ( .B0(n5000), .B1(n5532), .A0N(w_matrix[758]), .A1N(n5159), 
        .Y(n2677) );
  OAI2BB2X1 U6908 ( .B0(n5000), .B1(n5541), .A0N(w_matrix[822]), .A1N(n5168), 
        .Y(n2613) );
  OAI2BB2X1 U6909 ( .B0(n5000), .B1(n5576), .A0N(w_matrix[950]), .A1N(n5176), 
        .Y(n2485) );
  OAI2BB2X1 U6910 ( .B0(n4999), .B1(n5411), .A0N(w_matrix[55]), .A1N(n5096), 
        .Y(n3380) );
  OAI2BB2X1 U6911 ( .B0(n4999), .B1(n5433), .A0N(w_matrix[183]), .A1N(n5106), 
        .Y(n3252) );
  OAI2BB2X1 U6912 ( .B0(n4999), .B1(n5450), .A0N(w_matrix[311]), .A1N(n5116), 
        .Y(n3124) );
  OAI2BB2X1 U6913 ( .B0(n4999), .B1(n5463), .A0N(w_matrix[375]), .A1N(n5124), 
        .Y(n3060) );
  OAI2BB2X1 U6914 ( .B0(n4999), .B1(n5472), .A0N(w_matrix[439]), .A1N(n5132), 
        .Y(n2996) );
  OAI2BB2X1 U6915 ( .B0(n4999), .B1(n5485), .A0N(w_matrix[503]), .A1N(n5140), 
        .Y(n2932) );
  OAI2BB2X1 U6916 ( .B0(n4999), .B1(n5510), .A0N(w_matrix[631]), .A1N(n5148), 
        .Y(n2804) );
  OAI2BB2X1 U6917 ( .B0(n4999), .B1(n5532), .A0N(w_matrix[759]), .A1N(n5159), 
        .Y(n2676) );
  OAI2BB2X1 U6918 ( .B0(n4999), .B1(n5540), .A0N(w_matrix[823]), .A1N(n5168), 
        .Y(n2612) );
  OAI2BB2X1 U6919 ( .B0(n4999), .B1(n5575), .A0N(w_matrix[951]), .A1N(n5176), 
        .Y(n2484) );
  OAI2BB2X1 U6920 ( .B0(n4998), .B1(n5411), .A0N(w_matrix[56]), .A1N(n5096), 
        .Y(n3379) );
  OAI2BB2X1 U6921 ( .B0(n4998), .B1(n5433), .A0N(w_matrix[184]), .A1N(n5106), 
        .Y(n3251) );
  OAI2BB2X1 U6922 ( .B0(n4998), .B1(n5450), .A0N(w_matrix[312]), .A1N(n5116), 
        .Y(n3123) );
  OAI2BB2X1 U6923 ( .B0(n4998), .B1(n5472), .A0N(w_matrix[440]), .A1N(n5132), 
        .Y(n2995) );
  OAI2BB2X1 U6924 ( .B0(n4998), .B1(n5510), .A0N(w_matrix[632]), .A1N(n5148), 
        .Y(n2803) );
  OAI2BB2X1 U6925 ( .B0(n4998), .B1(n5532), .A0N(w_matrix[760]), .A1N(n5159), 
        .Y(n2675) );
  OAI2BB2X1 U6926 ( .B0(n4997), .B1(n5411), .A0N(w_matrix[57]), .A1N(n5096), 
        .Y(n3378) );
  OAI2BB2X1 U6927 ( .B0(n4997), .B1(n5433), .A0N(w_matrix[185]), .A1N(n5106), 
        .Y(n3250) );
  OAI2BB2X1 U6928 ( .B0(n4997), .B1(n5450), .A0N(w_matrix[313]), .A1N(n5116), 
        .Y(n3122) );
  OAI2BB2X1 U6929 ( .B0(n4997), .B1(n5472), .A0N(w_matrix[441]), .A1N(n5132), 
        .Y(n2994) );
  OAI2BB2X1 U6930 ( .B0(n4997), .B1(n5510), .A0N(w_matrix[633]), .A1N(n5148), 
        .Y(n2802) );
  OAI2BB2X1 U6931 ( .B0(n4997), .B1(n5532), .A0N(w_matrix[761]), .A1N(n5159), 
        .Y(n2674) );
  OAI2BB2X1 U6932 ( .B0(n4996), .B1(n5411), .A0N(w_matrix[58]), .A1N(n5096), 
        .Y(n3377) );
  OAI2BB2X1 U6933 ( .B0(n4996), .B1(n5433), .A0N(w_matrix[186]), .A1N(n5106), 
        .Y(n3249) );
  OAI2BB2X1 U6934 ( .B0(n4996), .B1(n5450), .A0N(w_matrix[314]), .A1N(n5116), 
        .Y(n3121) );
  OAI2BB2X1 U6935 ( .B0(n4996), .B1(n5472), .A0N(w_matrix[442]), .A1N(n5132), 
        .Y(n2993) );
  OAI2BB2X1 U6936 ( .B0(n4996), .B1(n5510), .A0N(w_matrix[634]), .A1N(n5148), 
        .Y(n2801) );
  OAI2BB2X1 U6937 ( .B0(n4996), .B1(n5532), .A0N(w_matrix[762]), .A1N(n5159), 
        .Y(n2673) );
  OAI2BB2X1 U6938 ( .B0(n4995), .B1(n5411), .A0N(w_matrix[59]), .A1N(n5096), 
        .Y(n3376) );
  OAI2BB2X1 U6939 ( .B0(n4995), .B1(n5433), .A0N(w_matrix[187]), .A1N(n5106), 
        .Y(n3248) );
  OAI2BB2X1 U6940 ( .B0(n4995), .B1(n5450), .A0N(w_matrix[315]), .A1N(n5116), 
        .Y(n3120) );
  OAI2BB2X1 U6941 ( .B0(n4995), .B1(n5472), .A0N(w_matrix[443]), .A1N(n5132), 
        .Y(n2992) );
  OAI2BB2X1 U6942 ( .B0(n4995), .B1(n5510), .A0N(w_matrix[635]), .A1N(n5148), 
        .Y(n2800) );
  OAI2BB2X1 U6943 ( .B0(n4995), .B1(n5532), .A0N(w_matrix[763]), .A1N(n5159), 
        .Y(n2672) );
  OAI2BB2X1 U6944 ( .B0(n4994), .B1(n5462), .A0N(w_matrix[325]), .A1N(n5120), 
        .Y(n3110) );
  OAI2BB2X1 U6945 ( .B0(n4994), .B1(n5484), .A0N(w_matrix[453]), .A1N(n5136), 
        .Y(n2982) );
  OAI2BB2X1 U6946 ( .B0(n4994), .B1(n5539), .A0N(w_matrix[773]), .A1N(n5164), 
        .Y(n2662) );
  OAI2BB2X1 U6947 ( .B0(n4994), .B1(n5574), .A0N(w_matrix[901]), .A1N(n5172), 
        .Y(n2534) );
  OAI2BB2X1 U6948 ( .B0(n4993), .B1(n5411), .A0N(w_matrix[60]), .A1N(n5096), 
        .Y(n3375) );
  OAI2BB2X1 U6949 ( .B0(n4993), .B1(n5433), .A0N(w_matrix[188]), .A1N(n5106), 
        .Y(n3247) );
  OAI2BB2X1 U6950 ( .B0(n4993), .B1(n5450), .A0N(w_matrix[316]), .A1N(n5116), 
        .Y(n3119) );
  OAI2BB2X1 U6951 ( .B0(n4993), .B1(n5472), .A0N(w_matrix[444]), .A1N(n5132), 
        .Y(n2991) );
  OAI2BB2X1 U6952 ( .B0(n4993), .B1(n5510), .A0N(w_matrix[636]), .A1N(n5148), 
        .Y(n2799) );
  OAI2BB2X1 U6953 ( .B0(n4993), .B1(n5532), .A0N(w_matrix[764]), .A1N(n5159), 
        .Y(n2671) );
  OAI2BB2X1 U6954 ( .B0(n4992), .B1(n5450), .A0N(w_matrix[317]), .A1N(n5116), 
        .Y(n3118) );
  OAI2BB2X1 U6955 ( .B0(n4992), .B1(n5472), .A0N(w_matrix[445]), .A1N(n5132), 
        .Y(n2990) );
  OAI2BB2X1 U6956 ( .B0(n4991), .B1(n5450), .A0N(w_matrix[318]), .A1N(n5116), 
        .Y(n3117) );
  OAI2BB2X1 U6957 ( .B0(n4991), .B1(n5472), .A0N(w_matrix[446]), .A1N(n5132), 
        .Y(n2989) );
  OAI2BB2X1 U6958 ( .B0(n4990), .B1(n5453), .A0N(w_matrix[319]), .A1N(n5116), 
        .Y(n3116) );
  OAI2BB2X1 U6959 ( .B0(n4990), .B1(n5461), .A0N(w_matrix[383]), .A1N(n5124), 
        .Y(n3052) );
  OAI2BB2X1 U6960 ( .B0(n4990), .B1(n5475), .A0N(w_matrix[447]), .A1N(n5132), 
        .Y(n2988) );
  OAI2BB2X1 U6961 ( .B0(n4990), .B1(n5483), .A0N(w_matrix[511]), .A1N(n5140), 
        .Y(n2924) );
  OAI2BB2X1 U6962 ( .B0(n4990), .B1(n5538), .A0N(w_matrix[831]), .A1N(n5168), 
        .Y(n2604) );
  OAI2BB2X1 U6963 ( .B0(n4990), .B1(n5573), .A0N(w_matrix[959]), .A1N(n5176), 
        .Y(n2476) );
  OAI2BB2X1 U6964 ( .B0(n4989), .B1(n5461), .A0N(w_matrix[326]), .A1N(n5120), 
        .Y(n3109) );
  OAI2BB2X1 U6965 ( .B0(n4989), .B1(n5483), .A0N(w_matrix[454]), .A1N(n5136), 
        .Y(n2981) );
  OAI2BB2X1 U6966 ( .B0(n4989), .B1(n5538), .A0N(w_matrix[774]), .A1N(n5164), 
        .Y(n2661) );
  OAI2BB2X1 U6967 ( .B0(n4989), .B1(n5573), .A0N(w_matrix[902]), .A1N(n5172), 
        .Y(n2533) );
  OAI2BB2X1 U6968 ( .B0(n4988), .B1(n5461), .A0N(w_matrix[327]), .A1N(n5120), 
        .Y(n3108) );
  OAI2BB2X1 U6969 ( .B0(n4988), .B1(n5483), .A0N(w_matrix[455]), .A1N(n5136), 
        .Y(n2980) );
  OAI2BB2X1 U6970 ( .B0(n4988), .B1(n5538), .A0N(w_matrix[775]), .A1N(n5164), 
        .Y(n2660) );
  OAI2BB2X1 U6971 ( .B0(n4988), .B1(n5573), .A0N(w_matrix[903]), .A1N(n5172), 
        .Y(n2532) );
  OAI2BB2X1 U6972 ( .B0(n4987), .B1(n5462), .A0N(w_matrix[328]), .A1N(n5120), 
        .Y(n3107) );
  OAI2BB2X1 U6973 ( .B0(n4987), .B1(n5484), .A0N(w_matrix[456]), .A1N(n5136), 
        .Y(n2979) );
  OAI2BB2X1 U6974 ( .B0(n4987), .B1(n5539), .A0N(w_matrix[776]), .A1N(n5164), 
        .Y(n2659) );
  OAI2BB2X1 U6975 ( .B0(n4987), .B1(n5574), .A0N(w_matrix[904]), .A1N(n5172), 
        .Y(n2531) );
  OAI2BB2X1 U6976 ( .B0(n4986), .B1(n5408), .A0N(w_matrix[9]), .A1N(n5093), 
        .Y(n3426) );
  OAI2BB2X1 U6977 ( .B0(n4986), .B1(n5430), .A0N(w_matrix[137]), .A1N(n5103), 
        .Y(n3298) );
  OAI2BB2X1 U6978 ( .B0(n4986), .B1(n5461), .A0N(w_matrix[329]), .A1N(n5120), 
        .Y(n3106) );
  OAI2BB2X1 U6979 ( .B0(n4986), .B1(n5483), .A0N(w_matrix[457]), .A1N(n5136), 
        .Y(n2978) );
  OAI2BB2X1 U6980 ( .B0(n4986), .B1(n5507), .A0N(w_matrix[585]), .A1N(n5145), 
        .Y(n2850) );
  OAI2BB2X1 U6981 ( .B0(n4986), .B1(n5526), .A0N(w_matrix[713]), .A1N(n5156), 
        .Y(n2722) );
  OAI2BB2X1 U6982 ( .B0(n4986), .B1(n5538), .A0N(w_matrix[777]), .A1N(n5164), 
        .Y(n2658) );
  OAI2BB2X1 U6983 ( .B0(n4986), .B1(n5573), .A0N(w_matrix[905]), .A1N(n5172), 
        .Y(n2530) );
  OAI2BB2X1 U6984 ( .B0(n5049), .B1(n5417), .A0N(w_matrix[64]), .A1N(n5342), 
        .Y(n3371) );
  OAI2BB2X1 U6985 ( .B0(n5049), .B1(n5439), .A0N(w_matrix[192]), .A1N(n5355), 
        .Y(n3243) );
  OAI2BB2X1 U6986 ( .B0(n5048), .B1(n5419), .A0N(w_matrix[74]), .A1N(n5339), 
        .Y(n3361) );
  OAI2BB2X1 U6987 ( .B0(n5048), .B1(n5441), .A0N(w_matrix[202]), .A1N(n5352), 
        .Y(n3233) );
  OAI2BB2X1 U6988 ( .B0(n5048), .B1(n5496), .A0N(w_matrix[522]), .A1N(n5363), 
        .Y(n2913) );
  OAI2BB2X1 U6989 ( .B0(n5048), .B1(n5518), .A0N(w_matrix[650]), .A1N(n5385), 
        .Y(n2785) );
  OAI2BB2X1 U6990 ( .B0(n5047), .B1(n5419), .A0N(w_matrix[75]), .A1N(n5340), 
        .Y(n3360) );
  OAI2BB2X1 U6991 ( .B0(n5047), .B1(n5441), .A0N(w_matrix[203]), .A1N(n5353), 
        .Y(n3232) );
  OAI2BB2X1 U6992 ( .B0(n5047), .B1(n5495), .A0N(w_matrix[523]), .A1N(n5363), 
        .Y(n2912) );
  OAI2BB2X1 U6993 ( .B0(n5047), .B1(n5517), .A0N(w_matrix[651]), .A1N(n5385), 
        .Y(n2784) );
  OAI2BB2X1 U6994 ( .B0(n5046), .B1(n5419), .A0N(w_matrix[76]), .A1N(n5344), 
        .Y(n3359) );
  OAI2BB2X1 U6995 ( .B0(n5046), .B1(n5441), .A0N(w_matrix[204]), .A1N(n5357), 
        .Y(n3231) );
  OAI2BB2X1 U6996 ( .B0(n5046), .B1(n5496), .A0N(w_matrix[524]), .A1N(n5363), 
        .Y(n2911) );
  OAI2BB2X1 U6997 ( .B0(n5046), .B1(n5518), .A0N(w_matrix[652]), .A1N(n5385), 
        .Y(n2783) );
  OAI2BB2X1 U6998 ( .B0(n5045), .B1(n5495), .A0N(w_matrix[525]), .A1N(n5363), 
        .Y(n2910) );
  OAI2BB2X1 U6999 ( .B0(n5045), .B1(n5517), .A0N(w_matrix[653]), .A1N(n5385), 
        .Y(n2782) );
  OAI2BB2X1 U7000 ( .B0(n5044), .B1(n5496), .A0N(w_matrix[526]), .A1N(n5363), 
        .Y(n2909) );
  OAI2BB2X1 U7001 ( .B0(n5044), .B1(n5518), .A0N(w_matrix[654]), .A1N(n5385), 
        .Y(n2781) );
  OAI2BB2X1 U7002 ( .B0(n5043), .B1(n5495), .A0N(w_matrix[527]), .A1N(n5363), 
        .Y(n2908) );
  OAI2BB2X1 U7003 ( .B0(n5043), .B1(n5517), .A0N(w_matrix[655]), .A1N(n5385), 
        .Y(n2780) );
  OAI2BB2X1 U7004 ( .B0(n5042), .B1(n5419), .A0N(w_matrix[80]), .A1N(n5344), 
        .Y(n3355) );
  OAI2BB2X1 U7005 ( .B0(n5042), .B1(n5441), .A0N(w_matrix[208]), .A1N(n5357), 
        .Y(n3227) );
  OAI2BB2X1 U7006 ( .B0(n5042), .B1(n5496), .A0N(w_matrix[528]), .A1N(n5363), 
        .Y(n2907) );
  OAI2BB2X1 U7007 ( .B0(n5042), .B1(n5518), .A0N(w_matrix[656]), .A1N(n5385), 
        .Y(n2779) );
  OAI2BB2X1 U7008 ( .B0(n5041), .B1(n5418), .A0N(w_matrix[81]), .A1N(n5341), 
        .Y(n3354) );
  OAI2BB2X1 U7009 ( .B0(n5041), .B1(n5440), .A0N(w_matrix[209]), .A1N(n5354), 
        .Y(n3226) );
  OAI2BB2X1 U7010 ( .B0(n5041), .B1(n5495), .A0N(w_matrix[529]), .A1N(n5363), 
        .Y(n2906) );
  OAI2BB2X1 U7011 ( .B0(n5041), .B1(n5517), .A0N(w_matrix[657]), .A1N(n5385), 
        .Y(n2778) );
  OAI2BB2X1 U7012 ( .B0(n5040), .B1(n5418), .A0N(w_matrix[82]), .A1N(n5341), 
        .Y(n3353) );
  OAI2BB2X1 U7013 ( .B0(n5040), .B1(n5440), .A0N(w_matrix[210]), .A1N(n5354), 
        .Y(n3225) );
  OAI2BB2X1 U7014 ( .B0(n5040), .B1(n5497), .A0N(w_matrix[530]), .A1N(n5364), 
        .Y(n2905) );
  OAI2BB2X1 U7015 ( .B0(n5040), .B1(n5519), .A0N(w_matrix[658]), .A1N(n5386), 
        .Y(n2777) );
  OAI2BB2X1 U7016 ( .B0(n5039), .B1(n5418), .A0N(w_matrix[83]), .A1N(n5341), 
        .Y(n3352) );
  OAI2BB2X1 U7017 ( .B0(n5039), .B1(n5440), .A0N(w_matrix[211]), .A1N(n5354), 
        .Y(n3224) );
  OAI2BB2X1 U7018 ( .B0(n5039), .B1(n5496), .A0N(w_matrix[531]), .A1N(n5364), 
        .Y(n2904) );
  OAI2BB2X1 U7019 ( .B0(n5039), .B1(n5518), .A0N(w_matrix[659]), .A1N(n5386), 
        .Y(n2776) );
  OAI2BB2X1 U7020 ( .B0(n5038), .B1(n5419), .A0N(w_matrix[65]), .A1N(n5339), 
        .Y(n3370) );
  OAI2BB2X1 U7021 ( .B0(n5038), .B1(n5441), .A0N(w_matrix[193]), .A1N(n5352), 
        .Y(n3242) );
  OAI2BB2X1 U7022 ( .B0(n5037), .B1(n5418), .A0N(w_matrix[84]), .A1N(n5341), 
        .Y(n3351) );
  OAI2BB2X1 U7023 ( .B0(n5037), .B1(n5440), .A0N(w_matrix[212]), .A1N(n5354), 
        .Y(n3223) );
  OAI2BB2X1 U7024 ( .B0(n5037), .B1(n5496), .A0N(w_matrix[532]), .A1N(n5364), 
        .Y(n2903) );
  OAI2BB2X1 U7025 ( .B0(n5037), .B1(n5518), .A0N(w_matrix[660]), .A1N(n5386), 
        .Y(n2775) );
  OAI2BB2X1 U7026 ( .B0(n5036), .B1(n5418), .A0N(w_matrix[85]), .A1N(n5345), 
        .Y(n3350) );
  OAI2BB2X1 U7027 ( .B0(n5036), .B1(n5440), .A0N(w_matrix[213]), .A1N(n5358), 
        .Y(n3222) );
  OAI2BB2X1 U7028 ( .B0(n5036), .B1(n5496), .A0N(w_matrix[533]), .A1N(n5364), 
        .Y(n2902) );
  OAI2BB2X1 U7029 ( .B0(n5036), .B1(n5518), .A0N(w_matrix[661]), .A1N(n5386), 
        .Y(n2774) );
  OAI2BB2X1 U7030 ( .B0(n5035), .B1(n5418), .A0N(w_matrix[86]), .A1N(n5346), 
        .Y(n3349) );
  OAI2BB2X1 U7031 ( .B0(n5035), .B1(n5440), .A0N(w_matrix[214]), .A1N(n5359), 
        .Y(n3221) );
  OAI2BB2X1 U7032 ( .B0(n5035), .B1(n5496), .A0N(w_matrix[534]), .A1N(n5364), 
        .Y(n2901) );
  OAI2BB2X1 U7033 ( .B0(n5035), .B1(n5518), .A0N(w_matrix[662]), .A1N(n5386), 
        .Y(n2773) );
  OAI2BB2X1 U7034 ( .B0(n5034), .B1(n5418), .A0N(w_matrix[87]), .A1N(n5339), 
        .Y(n3348) );
  OAI2BB2X1 U7035 ( .B0(n5034), .B1(n5440), .A0N(w_matrix[215]), .A1N(n5352), 
        .Y(n3220) );
  OAI2BB2X1 U7036 ( .B0(n5034), .B1(n5496), .A0N(w_matrix[535]), .A1N(n5364), 
        .Y(n2900) );
  OAI2BB2X1 U7037 ( .B0(n5034), .B1(n5518), .A0N(w_matrix[663]), .A1N(n5386), 
        .Y(n2772) );
  OAI2BB2X1 U7038 ( .B0(n5033), .B1(n5418), .A0N(w_matrix[88]), .A1N(n5340), 
        .Y(n3347) );
  OAI2BB2X1 U7039 ( .B0(n5033), .B1(n5440), .A0N(w_matrix[216]), .A1N(n5353), 
        .Y(n3219) );
  OAI2BB2X1 U7040 ( .B0(n5033), .B1(n5496), .A0N(w_matrix[536]), .A1N(n5364), 
        .Y(n2899) );
  OAI2BB2X1 U7041 ( .B0(n5033), .B1(n5518), .A0N(w_matrix[664]), .A1N(n5386), 
        .Y(n2771) );
  OAI2BB2X1 U7042 ( .B0(n5032), .B1(n5418), .A0N(w_matrix[89]), .A1N(n5342), 
        .Y(n3346) );
  OAI2BB2X1 U7043 ( .B0(n5032), .B1(n5440), .A0N(w_matrix[217]), .A1N(n5355), 
        .Y(n3218) );
  OAI2BB2X1 U7044 ( .B0(n5032), .B1(n5496), .A0N(w_matrix[537]), .A1N(n5364), 
        .Y(n2898) );
  OAI2BB2X1 U7045 ( .B0(n5032), .B1(n5518), .A0N(w_matrix[665]), .A1N(n5386), 
        .Y(n2770) );
  OAI2BB2X1 U7046 ( .B0(n5031), .B1(n5418), .A0N(w_matrix[90]), .A1N(n5342), 
        .Y(n3345) );
  OAI2BB2X1 U7047 ( .B0(n5031), .B1(n5440), .A0N(w_matrix[218]), .A1N(n5355), 
        .Y(n3217) );
  OAI2BB2X1 U7048 ( .B0(n5031), .B1(n5496), .A0N(w_matrix[538]), .A1N(n5364), 
        .Y(n2897) );
  OAI2BB2X1 U7049 ( .B0(n5031), .B1(n5518), .A0N(w_matrix[666]), .A1N(n5386), 
        .Y(n2769) );
  OAI2BB2X1 U7050 ( .B0(n5030), .B1(n5418), .A0N(w_matrix[91]), .A1N(n5342), 
        .Y(n3344) );
  OAI2BB2X1 U7051 ( .B0(n5030), .B1(n5440), .A0N(w_matrix[219]), .A1N(n5355), 
        .Y(n3216) );
  OAI2BB2X1 U7052 ( .B0(n5030), .B1(n5496), .A0N(w_matrix[539]), .A1N(n5364), 
        .Y(n2896) );
  OAI2BB2X1 U7053 ( .B0(n5030), .B1(n5518), .A0N(w_matrix[667]), .A1N(n5386), 
        .Y(n2768) );
  OAI2BB2X1 U7054 ( .B0(n5029), .B1(n5418), .A0N(w_matrix[92]), .A1N(n5342), 
        .Y(n3343) );
  OAI2BB2X1 U7055 ( .B0(n5029), .B1(n5440), .A0N(w_matrix[220]), .A1N(n5355), 
        .Y(n3215) );
  OAI2BB2X1 U7056 ( .B0(n5029), .B1(n5496), .A0N(w_matrix[540]), .A1N(n5364), 
        .Y(n2895) );
  OAI2BB2X1 U7057 ( .B0(n5029), .B1(n5518), .A0N(w_matrix[668]), .A1N(n5386), 
        .Y(n2767) );
  OAI2BB2X1 U7058 ( .B0(n5028), .B1(n5418), .A0N(w_matrix[93]), .A1N(n5340), 
        .Y(n3342) );
  OAI2BB2X1 U7059 ( .B0(n5028), .B1(n5440), .A0N(w_matrix[221]), .A1N(n5353), 
        .Y(n3214) );
  OAI2BB2X1 U7060 ( .B0(n5028), .B1(n5496), .A0N(w_matrix[541]), .A1N(n5364), 
        .Y(n2894) );
  OAI2BB2X1 U7061 ( .B0(n5028), .B1(n5518), .A0N(w_matrix[669]), .A1N(n5386), 
        .Y(n2766) );
  OAI2BB2X1 U7062 ( .B0(n5027), .B1(n5419), .A0N(w_matrix[66]), .A1N(n5339), 
        .Y(n3369) );
  OAI2BB2X1 U7063 ( .B0(n5027), .B1(n5441), .A0N(w_matrix[194]), .A1N(n5352), 
        .Y(n3241) );
  OAI2BB2X1 U7064 ( .B0(n5026), .B1(n5421), .A0N(w_matrix[94]), .A1N(n5342), 
        .Y(n3341) );
  OAI2BB2X1 U7065 ( .B0(n5026), .B1(n5443), .A0N(w_matrix[222]), .A1N(n5355), 
        .Y(n3213) );
  OAI2BB2X1 U7066 ( .B0(n5026), .B1(n5496), .A0N(w_matrix[542]), .A1N(n5364), 
        .Y(n2893) );
  OAI2BB2X1 U7067 ( .B0(n5026), .B1(n5518), .A0N(w_matrix[670]), .A1N(n5386), 
        .Y(n2765) );
  OAI2BB2X1 U7068 ( .B0(n5025), .B1(n5417), .A0N(w_matrix[95]), .A1N(n5345), 
        .Y(n3340) );
  OAI2BB2X1 U7069 ( .B0(n5025), .B1(n5439), .A0N(w_matrix[223]), .A1N(n5358), 
        .Y(n3212) );
  OAI2BB2X1 U7070 ( .B0(n5025), .B1(n5495), .A0N(w_matrix[543]), .A1N(n5365), 
        .Y(n2892) );
  OAI2BB2X1 U7071 ( .B0(n5025), .B1(n5517), .A0N(w_matrix[671]), .A1N(n5387), 
        .Y(n2764) );
  OAI2BB2X1 U7072 ( .B0(n5024), .B1(n5417), .A0N(w_matrix[96]), .A1N(n5339), 
        .Y(n3339) );
  OAI2BB2X1 U7073 ( .B0(n5024), .B1(n5439), .A0N(w_matrix[224]), .A1N(n5352), 
        .Y(n3211) );
  OAI2BB2X1 U7074 ( .B0(n5024), .B1(n5495), .A0N(w_matrix[544]), .A1N(n5365), 
        .Y(n2891) );
  OAI2BB2X1 U7075 ( .B0(n5024), .B1(n5517), .A0N(w_matrix[672]), .A1N(n5387), 
        .Y(n2763) );
  OAI2BB2X1 U7076 ( .B0(n5023), .B1(n5421), .A0N(w_matrix[97]), .A1N(n5343), 
        .Y(n3338) );
  OAI2BB2X1 U7077 ( .B0(n5023), .B1(n5443), .A0N(w_matrix[225]), .A1N(n5356), 
        .Y(n3210) );
  OAI2BB2X1 U7078 ( .B0(n5023), .B1(n5495), .A0N(w_matrix[545]), .A1N(n5365), 
        .Y(n2890) );
  OAI2BB2X1 U7079 ( .B0(n5023), .B1(n5517), .A0N(w_matrix[673]), .A1N(n5387), 
        .Y(n2762) );
  OAI2BB2X1 U7080 ( .B0(n5022), .B1(n5417), .A0N(w_matrix[98]), .A1N(n5343), 
        .Y(n3337) );
  OAI2BB2X1 U7081 ( .B0(n5022), .B1(n5439), .A0N(w_matrix[226]), .A1N(n5356), 
        .Y(n3209) );
  OAI2BB2X1 U7082 ( .B0(n5022), .B1(n5495), .A0N(w_matrix[546]), .A1N(n5365), 
        .Y(n2889) );
  OAI2BB2X1 U7083 ( .B0(n5022), .B1(n5517), .A0N(w_matrix[674]), .A1N(n5387), 
        .Y(n2761) );
  OAI2BB2X1 U7084 ( .B0(n5021), .B1(n5421), .A0N(w_matrix[99]), .A1N(n5343), 
        .Y(n3336) );
  OAI2BB2X1 U7085 ( .B0(n5021), .B1(n5443), .A0N(w_matrix[227]), .A1N(n5356), 
        .Y(n3208) );
  OAI2BB2X1 U7086 ( .B0(n5021), .B1(n5495), .A0N(w_matrix[547]), .A1N(n5365), 
        .Y(n2888) );
  OAI2BB2X1 U7087 ( .B0(n5021), .B1(n5517), .A0N(w_matrix[675]), .A1N(n5387), 
        .Y(n2760) );
  OAI2BB2X1 U7088 ( .B0(n5020), .B1(n5417), .A0N(w_matrix[100]), .A1N(n5343), 
        .Y(n3335) );
  OAI2BB2X1 U7089 ( .B0(n5020), .B1(n5439), .A0N(w_matrix[228]), .A1N(n5356), 
        .Y(n3207) );
  OAI2BB2X1 U7090 ( .B0(n5020), .B1(n5495), .A0N(w_matrix[548]), .A1N(n5365), 
        .Y(n2887) );
  OAI2BB2X1 U7091 ( .B0(n5020), .B1(n5517), .A0N(w_matrix[676]), .A1N(n5387), 
        .Y(n2759) );
  OAI2BB2X1 U7092 ( .B0(n5019), .B1(n5420), .A0N(w_matrix[101]), .A1N(n5344), 
        .Y(n3334) );
  OAI2BB2X1 U7093 ( .B0(n5019), .B1(n5442), .A0N(w_matrix[229]), .A1N(n5357), 
        .Y(n3206) );
  OAI2BB2X1 U7094 ( .B0(n5019), .B1(n5494), .A0N(w_matrix[549]), .A1N(n5365), 
        .Y(n2886) );
  OAI2BB2X1 U7095 ( .B0(n5019), .B1(n5516), .A0N(w_matrix[677]), .A1N(n5387), 
        .Y(n2758) );
  OAI2BB2X1 U7096 ( .B0(n5018), .B1(n5418), .A0N(w_matrix[102]), .A1N(n5344), 
        .Y(n3333) );
  OAI2BB2X1 U7097 ( .B0(n5018), .B1(n5440), .A0N(w_matrix[230]), .A1N(n5357), 
        .Y(n3205) );
  OAI2BB2X1 U7098 ( .B0(n5018), .B1(n5495), .A0N(w_matrix[550]), .A1N(n5365), 
        .Y(n2885) );
  OAI2BB2X1 U7099 ( .B0(n5018), .B1(n5517), .A0N(w_matrix[678]), .A1N(n5387), 
        .Y(n2757) );
  OAI2BB2X1 U7100 ( .B0(n5017), .B1(n5419), .A0N(w_matrix[103]), .A1N(n5344), 
        .Y(n3332) );
  OAI2BB2X1 U7101 ( .B0(n5017), .B1(n5441), .A0N(w_matrix[231]), .A1N(n5357), 
        .Y(n3204) );
  OAI2BB2X1 U7102 ( .B0(n5017), .B1(n5494), .A0N(w_matrix[551]), .A1N(n5365), 
        .Y(n2884) );
  OAI2BB2X1 U7103 ( .B0(n5017), .B1(n5516), .A0N(w_matrix[679]), .A1N(n5387), 
        .Y(n2756) );
  OAI2BB2X1 U7104 ( .B0(n5016), .B1(n5419), .A0N(w_matrix[67]), .A1N(n5339), 
        .Y(n3368) );
  OAI2BB2X1 U7105 ( .B0(n5016), .B1(n5441), .A0N(w_matrix[195]), .A1N(n5352), 
        .Y(n3240) );
  OAI2BB2X1 U7106 ( .B0(n5015), .B1(n5416), .A0N(w_matrix[104]), .A1N(n5344), 
        .Y(n3331) );
  OAI2BB2X1 U7107 ( .B0(n5015), .B1(n5438), .A0N(w_matrix[232]), .A1N(n5357), 
        .Y(n3203) );
  OAI2BB2X1 U7108 ( .B0(n5015), .B1(n5495), .A0N(w_matrix[552]), .A1N(n5365), 
        .Y(n2883) );
  OAI2BB2X1 U7109 ( .B0(n5015), .B1(n5517), .A0N(w_matrix[680]), .A1N(n5387), 
        .Y(n2755) );
  OAI2BB2X1 U7110 ( .B0(n5014), .B1(n5420), .A0N(w_matrix[105]), .A1N(n5345), 
        .Y(n3330) );
  OAI2BB2X1 U7111 ( .B0(n5014), .B1(n5442), .A0N(w_matrix[233]), .A1N(n5358), 
        .Y(n3202) );
  OAI2BB2X1 U7112 ( .B0(n5014), .B1(n5494), .A0N(w_matrix[553]), .A1N(n5365), 
        .Y(n2882) );
  OAI2BB2X1 U7113 ( .B0(n5014), .B1(n5516), .A0N(w_matrix[681]), .A1N(n5387), 
        .Y(n2754) );
  OAI2BB2X1 U7114 ( .B0(n5013), .B1(n5415), .A0N(w_matrix[106]), .A1N(n5345), 
        .Y(n3329) );
  OAI2BB2X1 U7115 ( .B0(n5013), .B1(n5437), .A0N(w_matrix[234]), .A1N(n5358), 
        .Y(n3201) );
  OAI2BB2X1 U7116 ( .B0(n5013), .B1(n5495), .A0N(w_matrix[554]), .A1N(n5365), 
        .Y(n2881) );
  OAI2BB2X1 U7117 ( .B0(n5013), .B1(n5517), .A0N(w_matrix[682]), .A1N(n5387), 
        .Y(n2753) );
  OAI2BB2X1 U7118 ( .B0(n5012), .B1(n5417), .A0N(w_matrix[107]), .A1N(n5345), 
        .Y(n3328) );
  OAI2BB2X1 U7119 ( .B0(n5012), .B1(n5439), .A0N(w_matrix[235]), .A1N(n5358), 
        .Y(n3200) );
  OAI2BB2X1 U7120 ( .B0(n5012), .B1(n5494), .A0N(w_matrix[555]), .A1N(n5365), 
        .Y(n2880) );
  OAI2BB2X1 U7121 ( .B0(n5012), .B1(n5516), .A0N(w_matrix[683]), .A1N(n5387), 
        .Y(n2752) );
  OAI2BB2X1 U7122 ( .B0(n5011), .B1(n5417), .A0N(w_matrix[108]), .A1N(n5345), 
        .Y(n3327) );
  OAI2BB2X1 U7123 ( .B0(n5011), .B1(n5439), .A0N(w_matrix[236]), .A1N(n5358), 
        .Y(n3199) );
  OAI2BB2X1 U7124 ( .B0(n5011), .B1(n5495), .A0N(w_matrix[556]), .A1N(n5366), 
        .Y(n2879) );
  OAI2BB2X1 U7125 ( .B0(n5011), .B1(n5517), .A0N(w_matrix[684]), .A1N(n5388), 
        .Y(n2751) );
  OAI2BB2X1 U7126 ( .B0(n5010), .B1(n5417), .A0N(w_matrix[109]), .A1N(n5346), 
        .Y(n3326) );
  OAI2BB2X1 U7127 ( .B0(n5010), .B1(n5439), .A0N(w_matrix[237]), .A1N(n5359), 
        .Y(n3198) );
  OAI2BB2X1 U7128 ( .B0(n5010), .B1(n5496), .A0N(w_matrix[557]), .A1N(n5366), 
        .Y(n2878) );
  OAI2BB2X1 U7129 ( .B0(n5010), .B1(n5518), .A0N(w_matrix[685]), .A1N(n5388), 
        .Y(n2750) );
  OAI2BB2X1 U7130 ( .B0(n5009), .B1(n5417), .A0N(w_matrix[110]), .A1N(n5346), 
        .Y(n3325) );
  OAI2BB2X1 U7131 ( .B0(n5009), .B1(n5439), .A0N(w_matrix[238]), .A1N(n5359), 
        .Y(n3197) );
  OAI2BB2X1 U7132 ( .B0(n5009), .B1(n5494), .A0N(w_matrix[558]), .A1N(n5366), 
        .Y(n2877) );
  OAI2BB2X1 U7133 ( .B0(n5009), .B1(n5516), .A0N(w_matrix[686]), .A1N(n5388), 
        .Y(n2749) );
  OAI2BB2X1 U7134 ( .B0(n5008), .B1(n5417), .A0N(w_matrix[111]), .A1N(n5346), 
        .Y(n3324) );
  OAI2BB2X1 U7135 ( .B0(n5008), .B1(n5439), .A0N(w_matrix[239]), .A1N(n5359), 
        .Y(n3196) );
  OAI2BB2X1 U7136 ( .B0(n5008), .B1(n5494), .A0N(w_matrix[559]), .A1N(n5366), 
        .Y(n2876) );
  OAI2BB2X1 U7137 ( .B0(n5008), .B1(n5516), .A0N(w_matrix[687]), .A1N(n5388), 
        .Y(n2748) );
  OAI2BB2X1 U7138 ( .B0(n5007), .B1(n5417), .A0N(w_matrix[112]), .A1N(n5346), 
        .Y(n3323) );
  OAI2BB2X1 U7139 ( .B0(n5007), .B1(n5439), .A0N(w_matrix[240]), .A1N(n5359), 
        .Y(n3195) );
  OAI2BB2X1 U7140 ( .B0(n5007), .B1(n5495), .A0N(w_matrix[560]), .A1N(n5366), 
        .Y(n2875) );
  OAI2BB2X1 U7141 ( .B0(n5007), .B1(n5517), .A0N(w_matrix[688]), .A1N(n5388), 
        .Y(n2747) );
  OAI2BB2X1 U7142 ( .B0(n5006), .B1(n5417), .A0N(w_matrix[113]), .A1N(n5341), 
        .Y(n3322) );
  OAI2BB2X1 U7143 ( .B0(n5006), .B1(n5439), .A0N(w_matrix[241]), .A1N(n5354), 
        .Y(n3194) );
  OAI2BB2X1 U7144 ( .B0(n5006), .B1(n5494), .A0N(w_matrix[561]), .A1N(n5366), 
        .Y(n2874) );
  OAI2BB2X1 U7145 ( .B0(n5006), .B1(n5516), .A0N(w_matrix[689]), .A1N(n5388), 
        .Y(n2746) );
  OAI2BB2X1 U7146 ( .B0(n5005), .B1(n5419), .A0N(w_matrix[68]), .A1N(n5339), 
        .Y(n3367) );
  OAI2BB2X1 U7147 ( .B0(n5005), .B1(n5441), .A0N(w_matrix[196]), .A1N(n5352), 
        .Y(n3239) );
  OAI2BB2X1 U7148 ( .B0(n5004), .B1(n5417), .A0N(w_matrix[114]), .A1N(n5337), 
        .Y(n3321) );
  OAI2BB2X1 U7149 ( .B0(n5004), .B1(n5439), .A0N(w_matrix[242]), .A1N(n5350), 
        .Y(n3193) );
  OAI2BB2X1 U7150 ( .B0(n5004), .B1(n5494), .A0N(w_matrix[562]), .A1N(n5366), 
        .Y(n2873) );
  OAI2BB2X1 U7151 ( .B0(n5004), .B1(n5516), .A0N(w_matrix[690]), .A1N(n5388), 
        .Y(n2745) );
  OAI2BB2X1 U7152 ( .B0(n5003), .B1(n5417), .A0N(w_matrix[115]), .A1N(n5342), 
        .Y(n3320) );
  OAI2BB2X1 U7153 ( .B0(n5003), .B1(n5439), .A0N(w_matrix[243]), .A1N(n5355), 
        .Y(n3192) );
  OAI2BB2X1 U7154 ( .B0(n5003), .B1(n5494), .A0N(w_matrix[563]), .A1N(n5366), 
        .Y(n2872) );
  OAI2BB2X1 U7155 ( .B0(n5003), .B1(n5516), .A0N(w_matrix[691]), .A1N(n5388), 
        .Y(n2744) );
  OAI2BB2X1 U7156 ( .B0(n5002), .B1(n5417), .A0N(w_matrix[116]), .A1N(n5339), 
        .Y(n3319) );
  OAI2BB2X1 U7157 ( .B0(n5002), .B1(n5439), .A0N(w_matrix[244]), .A1N(n5352), 
        .Y(n3191) );
  OAI2BB2X1 U7158 ( .B0(n5002), .B1(n5494), .A0N(w_matrix[564]), .A1N(n5366), 
        .Y(n2871) );
  OAI2BB2X1 U7159 ( .B0(n5002), .B1(n5516), .A0N(w_matrix[692]), .A1N(n5388), 
        .Y(n2743) );
  OAI2BB2X1 U7160 ( .B0(n5001), .B1(n5417), .A0N(w_matrix[117]), .A1N(n5340), 
        .Y(n3318) );
  OAI2BB2X1 U7161 ( .B0(n5001), .B1(n5439), .A0N(w_matrix[245]), .A1N(n5353), 
        .Y(n3190) );
  OAI2BB2X1 U7162 ( .B0(n5000), .B1(n5417), .A0N(w_matrix[118]), .A1N(n5345), 
        .Y(n3317) );
  OAI2BB2X1 U7163 ( .B0(n5000), .B1(n5439), .A0N(w_matrix[246]), .A1N(n5358), 
        .Y(n3189) );
  OAI2BB2X1 U7164 ( .B0(n5000), .B1(n5495), .A0N(w_matrix[566]), .A1N(n5366), 
        .Y(n2869) );
  OAI2BB2X1 U7165 ( .B0(n5000), .B1(n5517), .A0N(w_matrix[694]), .A1N(n5388), 
        .Y(n2741) );
  OAI2BB2X1 U7166 ( .B0(n4998), .B1(n5494), .A0N(w_matrix[568]), .A1N(n5366), 
        .Y(n2867) );
  OAI2BB2X1 U7167 ( .B0(n4998), .B1(n5516), .A0N(w_matrix[696]), .A1N(n5388), 
        .Y(n2739) );
  OAI2BB2X1 U7168 ( .B0(n4996), .B1(n5494), .A0N(w_matrix[570]), .A1N(n5367), 
        .Y(n2865) );
  OAI2BB2X1 U7169 ( .B0(n4996), .B1(n5516), .A0N(w_matrix[698]), .A1N(n5389), 
        .Y(n2737) );
  OAI2BB2X1 U7170 ( .B0(n4994), .B1(n5419), .A0N(w_matrix[69]), .A1N(n5340), 
        .Y(n3366) );
  OAI2BB2X1 U7171 ( .B0(n4994), .B1(n5441), .A0N(w_matrix[197]), .A1N(n5353), 
        .Y(n3238) );
  OAI2BB2X1 U7172 ( .B0(n4993), .B1(n5495), .A0N(w_matrix[572]), .A1N(n5367), 
        .Y(n2863) );
  OAI2BB2X1 U7173 ( .B0(n4993), .B1(n5517), .A0N(w_matrix[700]), .A1N(n5389), 
        .Y(n2735) );
  OAI2BB2X1 U7174 ( .B0(n4991), .B1(n5494), .A0N(w_matrix[574]), .A1N(n5367), 
        .Y(n2861) );
  OAI2BB2X1 U7175 ( .B0(n4991), .B1(n5516), .A0N(w_matrix[702]), .A1N(n5389), 
        .Y(n2733) );
  OAI2BB2X1 U7176 ( .B0(n4990), .B1(n5499), .A0N(w_matrix[575]), .A1N(n5367), 
        .Y(n2860) );
  OAI2BB2X1 U7177 ( .B0(n4990), .B1(n5521), .A0N(w_matrix[703]), .A1N(n5389), 
        .Y(n2732) );
  OAI2BB2X1 U7178 ( .B0(n4989), .B1(n5419), .A0N(w_matrix[70]), .A1N(n5340), 
        .Y(n3365) );
  OAI2BB2X1 U7179 ( .B0(n4989), .B1(n5441), .A0N(w_matrix[198]), .A1N(n5353), 
        .Y(n3237) );
  OAI2BB2X1 U7180 ( .B0(n4988), .B1(n5419), .A0N(w_matrix[71]), .A1N(n5340), 
        .Y(n3364) );
  OAI2BB2X1 U7181 ( .B0(n4988), .B1(n5441), .A0N(w_matrix[199]), .A1N(n5353), 
        .Y(n3236) );
  OAI2BB2X1 U7182 ( .B0(n4988), .B1(n5498), .A0N(w_matrix[519]), .A1N(n5363), 
        .Y(n2916) );
  OAI2BB2X1 U7183 ( .B0(n4988), .B1(n5520), .A0N(w_matrix[647]), .A1N(n5385), 
        .Y(n2788) );
  OAI2BB2X1 U7184 ( .B0(n4987), .B1(n5419), .A0N(w_matrix[72]), .A1N(n5340), 
        .Y(n3363) );
  OAI2BB2X1 U7185 ( .B0(n4987), .B1(n5441), .A0N(w_matrix[200]), .A1N(n5353), 
        .Y(n3235) );
  OAI2BB2X1 U7186 ( .B0(n4987), .B1(n5497), .A0N(w_matrix[520]), .A1N(n5363), 
        .Y(n2915) );
  OAI2BB2X1 U7187 ( .B0(n4987), .B1(n5519), .A0N(w_matrix[648]), .A1N(n5385), 
        .Y(n2787) );
  OAI2BB2X1 U7188 ( .B0(n4986), .B1(n5419), .A0N(w_matrix[73]), .A1N(n5346), 
        .Y(n3362) );
  OAI2BB2X1 U7189 ( .B0(n4986), .B1(n5441), .A0N(w_matrix[201]), .A1N(n5359), 
        .Y(n3234) );
  OAI2BB2X1 U7190 ( .B0(n4986), .B1(n5492), .A0N(w_matrix[521]), .A1N(n5363), 
        .Y(n2914) );
  OAI2BB2X1 U7191 ( .B0(n4986), .B1(n5514), .A0N(w_matrix[649]), .A1N(n5385), 
        .Y(n2786) );
  OAI2BB2X1 U7192 ( .B0(n5049), .B1(n5454), .A0N(w_matrix[256]), .A1N(n5112), 
        .Y(n3179) );
  OAI2BB2X1 U7193 ( .B0(n5049), .B1(n5476), .A0N(w_matrix[384]), .A1N(n5128), 
        .Y(n3051) );
  OAI2BB2X1 U7194 ( .B0(n5048), .B1(n5454), .A0N(w_matrix[266]), .A1N(n5112), 
        .Y(n3169) );
  OAI2BB2X1 U7195 ( .B0(n5048), .B1(n5476), .A0N(w_matrix[394]), .A1N(n5128), 
        .Y(n3041) );
  OAI2BB2X1 U7196 ( .B0(n5047), .B1(n5454), .A0N(w_matrix[267]), .A1N(n5112), 
        .Y(n3168) );
  OAI2BB2X1 U7197 ( .B0(n5047), .B1(n5476), .A0N(w_matrix[395]), .A1N(n5128), 
        .Y(n3040) );
  OAI2BB2X1 U7198 ( .B0(n5038), .B1(n5454), .A0N(w_matrix[257]), .A1N(n5112), 
        .Y(n3178) );
  OAI2BB2X1 U7199 ( .B0(n5038), .B1(n5476), .A0N(w_matrix[385]), .A1N(n5128), 
        .Y(n3050) );
  OAI2BB2X1 U7200 ( .B0(n5027), .B1(n5454), .A0N(w_matrix[258]), .A1N(n5112), 
        .Y(n3177) );
  OAI2BB2X1 U7201 ( .B0(n5027), .B1(n5476), .A0N(w_matrix[386]), .A1N(n5128), 
        .Y(n3049) );
  OAI2BB2X1 U7202 ( .B0(n5016), .B1(n5454), .A0N(w_matrix[259]), .A1N(n5112), 
        .Y(n3176) );
  OAI2BB2X1 U7203 ( .B0(n5016), .B1(n5476), .A0N(w_matrix[387]), .A1N(n5128), 
        .Y(n3048) );
  OAI2BB2X1 U7204 ( .B0(n5009), .B1(n5465), .A0N(w_matrix[366]), .A1N(n5123), 
        .Y(n3069) );
  OAI2BB2X1 U7205 ( .B0(n5009), .B1(n5487), .A0N(w_matrix[494]), .A1N(n5139), 
        .Y(n2941) );
  OAI2BB2X1 U7206 ( .B0(n5009), .B1(n5542), .A0N(w_matrix[814]), .A1N(n5167), 
        .Y(n2621) );
  OAI2BB2X1 U7207 ( .B0(n5009), .B1(n5577), .A0N(w_matrix[942]), .A1N(n5175), 
        .Y(n2493) );
  OAI2BB2X1 U7208 ( .B0(n5006), .B1(n5465), .A0N(w_matrix[369]), .A1N(n5123), 
        .Y(n3066) );
  OAI2BB2X1 U7209 ( .B0(n5006), .B1(n5487), .A0N(w_matrix[497]), .A1N(n5139), 
        .Y(n2938) );
  OAI2BB2X1 U7210 ( .B0(n5006), .B1(n5542), .A0N(w_matrix[817]), .A1N(n5167), 
        .Y(n2618) );
  OAI2BB2X1 U7211 ( .B0(n5006), .B1(n5577), .A0N(w_matrix[945]), .A1N(n5175), 
        .Y(n2490) );
  OAI2BB2X1 U7212 ( .B0(n5005), .B1(n5454), .A0N(w_matrix[260]), .A1N(n5112), 
        .Y(n3175) );
  OAI2BB2X1 U7213 ( .B0(n5005), .B1(n5476), .A0N(w_matrix[388]), .A1N(n5128), 
        .Y(n3047) );
  OAI2BB2X1 U7214 ( .B0(n5004), .B1(n5465), .A0N(w_matrix[370]), .A1N(n5123), 
        .Y(n3065) );
  OAI2BB2X1 U7215 ( .B0(n5004), .B1(n5487), .A0N(w_matrix[498]), .A1N(n5139), 
        .Y(n2937) );
  OAI2BB2X1 U7216 ( .B0(n5004), .B1(n5542), .A0N(w_matrix[818]), .A1N(n5167), 
        .Y(n2617) );
  OAI2BB2X1 U7217 ( .B0(n5004), .B1(n5577), .A0N(w_matrix[946]), .A1N(n5175), 
        .Y(n2489) );
  OAI2BB2X1 U7218 ( .B0(n5002), .B1(n5465), .A0N(w_matrix[372]), .A1N(n5124), 
        .Y(n3063) );
  OAI2BB2X1 U7219 ( .B0(n5002), .B1(n5487), .A0N(w_matrix[500]), .A1N(n5140), 
        .Y(n2935) );
  OAI2BB2X1 U7220 ( .B0(n5002), .B1(n5542), .A0N(w_matrix[820]), .A1N(n5168), 
        .Y(n2615) );
  OAI2BB2X1 U7221 ( .B0(n5002), .B1(n5577), .A0N(w_matrix[948]), .A1N(n5176), 
        .Y(n2487) );
  OAI2BB2X1 U7222 ( .B0(n5001), .B1(n5465), .A0N(w_matrix[373]), .A1N(n5124), 
        .Y(n3062) );
  OAI2BB2X1 U7223 ( .B0(n5001), .B1(n5487), .A0N(w_matrix[501]), .A1N(n5140), 
        .Y(n2934) );
  OAI2BB2X1 U7224 ( .B0(n5001), .B1(n5542), .A0N(w_matrix[821]), .A1N(n5168), 
        .Y(n2614) );
  OAI2BB2X1 U7225 ( .B0(n5001), .B1(n5577), .A0N(w_matrix[949]), .A1N(n5176), 
        .Y(n2486) );
  OAI2BB2X1 U7226 ( .B0(n4998), .B1(n5465), .A0N(w_matrix[376]), .A1N(n5124), 
        .Y(n3059) );
  OAI2BB2X1 U7227 ( .B0(n4998), .B1(n5487), .A0N(w_matrix[504]), .A1N(n5140), 
        .Y(n2931) );
  OAI2BB2X1 U7228 ( .B0(n4998), .B1(n5542), .A0N(w_matrix[824]), .A1N(n5168), 
        .Y(n2611) );
  OAI2BB2X1 U7229 ( .B0(n4998), .B1(n5577), .A0N(w_matrix[952]), .A1N(n5176), 
        .Y(n2483) );
  OAI2BB2X1 U7230 ( .B0(n4997), .B1(n5465), .A0N(w_matrix[377]), .A1N(n5124), 
        .Y(n3058) );
  OAI2BB2X1 U7231 ( .B0(n4997), .B1(n5487), .A0N(w_matrix[505]), .A1N(n5140), 
        .Y(n2930) );
  OAI2BB2X1 U7232 ( .B0(n4997), .B1(n5542), .A0N(w_matrix[825]), .A1N(n5168), 
        .Y(n2610) );
  OAI2BB2X1 U7233 ( .B0(n4997), .B1(n5577), .A0N(w_matrix[953]), .A1N(n5176), 
        .Y(n2482) );
  OAI2BB2X1 U7234 ( .B0(n4996), .B1(n5465), .A0N(w_matrix[378]), .A1N(n5124), 
        .Y(n3057) );
  OAI2BB2X1 U7235 ( .B0(n4996), .B1(n5487), .A0N(w_matrix[506]), .A1N(n5140), 
        .Y(n2929) );
  OAI2BB2X1 U7236 ( .B0(n4996), .B1(n5542), .A0N(w_matrix[826]), .A1N(n5168), 
        .Y(n2609) );
  OAI2BB2X1 U7237 ( .B0(n4996), .B1(n5577), .A0N(w_matrix[954]), .A1N(n5176), 
        .Y(n2481) );
  OAI2BB2X1 U7238 ( .B0(n4995), .B1(n5465), .A0N(w_matrix[379]), .A1N(n5124), 
        .Y(n3056) );
  OAI2BB2X1 U7239 ( .B0(n4995), .B1(n5487), .A0N(w_matrix[507]), .A1N(n5140), 
        .Y(n2928) );
  OAI2BB2X1 U7240 ( .B0(n4995), .B1(n5542), .A0N(w_matrix[827]), .A1N(n5168), 
        .Y(n2608) );
  OAI2BB2X1 U7241 ( .B0(n4995), .B1(n5577), .A0N(w_matrix[955]), .A1N(n5176), 
        .Y(n2480) );
  OAI2BB2X1 U7242 ( .B0(n4994), .B1(n5454), .A0N(w_matrix[261]), .A1N(n5112), 
        .Y(n3174) );
  OAI2BB2X1 U7243 ( .B0(n4994), .B1(n5476), .A0N(w_matrix[389]), .A1N(n5128), 
        .Y(n3046) );
  OAI2BB2X1 U7244 ( .B0(n4993), .B1(n5465), .A0N(w_matrix[380]), .A1N(n5124), 
        .Y(n3055) );
  OAI2BB2X1 U7245 ( .B0(n4993), .B1(n5487), .A0N(w_matrix[508]), .A1N(n5140), 
        .Y(n2927) );
  OAI2BB2X1 U7246 ( .B0(n4993), .B1(n5542), .A0N(w_matrix[828]), .A1N(n5168), 
        .Y(n2607) );
  OAI2BB2X1 U7247 ( .B0(n4993), .B1(n5577), .A0N(w_matrix[956]), .A1N(n5176), 
        .Y(n2479) );
  OAI2BB2X1 U7248 ( .B0(n4992), .B1(n5465), .A0N(w_matrix[381]), .A1N(n5124), 
        .Y(n3054) );
  OAI2BB2X1 U7249 ( .B0(n4992), .B1(n5487), .A0N(w_matrix[509]), .A1N(n5140), 
        .Y(n2926) );
  OAI2BB2X1 U7250 ( .B0(n4992), .B1(n5542), .A0N(w_matrix[829]), .A1N(n5168), 
        .Y(n2606) );
  OAI2BB2X1 U7251 ( .B0(n4992), .B1(n5577), .A0N(w_matrix[957]), .A1N(n5176), 
        .Y(n2478) );
  OAI2BB2X1 U7252 ( .B0(n4991), .B1(n5465), .A0N(w_matrix[382]), .A1N(n5124), 
        .Y(n3053) );
  OAI2BB2X1 U7253 ( .B0(n4991), .B1(n5487), .A0N(w_matrix[510]), .A1N(n5140), 
        .Y(n2925) );
  OAI2BB2X1 U7254 ( .B0(n4991), .B1(n5542), .A0N(w_matrix[830]), .A1N(n5168), 
        .Y(n2605) );
  OAI2BB2X1 U7255 ( .B0(n4991), .B1(n5577), .A0N(w_matrix[958]), .A1N(n5176), 
        .Y(n2477) );
  OAI2BB2X1 U7256 ( .B0(n4989), .B1(n5454), .A0N(w_matrix[262]), .A1N(n5112), 
        .Y(n3173) );
  OAI2BB2X1 U7257 ( .B0(n4989), .B1(n5476), .A0N(w_matrix[390]), .A1N(n5128), 
        .Y(n3045) );
  OAI2BB2X1 U7258 ( .B0(n4988), .B1(n5454), .A0N(w_matrix[263]), .A1N(n5112), 
        .Y(n3172) );
  OAI2BB2X1 U7259 ( .B0(n4988), .B1(n5476), .A0N(w_matrix[391]), .A1N(n5128), 
        .Y(n3044) );
  OAI2BB2X1 U7260 ( .B0(n4987), .B1(n5454), .A0N(w_matrix[264]), .A1N(n5112), 
        .Y(n3171) );
  OAI2BB2X1 U7261 ( .B0(n4987), .B1(n5476), .A0N(w_matrix[392]), .A1N(n5128), 
        .Y(n3043) );
  OAI2BB2X1 U7262 ( .B0(n4986), .B1(n5454), .A0N(w_matrix[265]), .A1N(n5112), 
        .Y(n3170) );
  OAI2BB2X1 U7263 ( .B0(n4986), .B1(n5476), .A0N(w_matrix[393]), .A1N(n5128), 
        .Y(n3042) );
  OAI2BB2X1 U7264 ( .B0(n5049), .B1(n5407), .A0N(w_matrix[0]), .A1N(n5092), 
        .Y(n3435) );
  OAI2BB2X1 U7265 ( .B0(n5049), .B1(n5429), .A0N(w_matrix[128]), .A1N(n5102), 
        .Y(n3307) );
  OAI2BB2X1 U7266 ( .B0(n5049), .B1(n5506), .A0N(w_matrix[576]), .A1N(n5144), 
        .Y(n2859) );
  OAI2BB2X1 U7267 ( .B0(n5049), .B1(n5529), .A0N(w_matrix[704]), .A1N(n5155), 
        .Y(n2731) );
  OAI2BB2X1 U7268 ( .B0(n5038), .B1(n5407), .A0N(w_matrix[1]), .A1N(n5092), 
        .Y(n3434) );
  OAI2BB2X1 U7269 ( .B0(n5038), .B1(n5429), .A0N(w_matrix[129]), .A1N(n5102), 
        .Y(n3306) );
  OAI2BB2X1 U7270 ( .B0(n5038), .B1(n5506), .A0N(w_matrix[577]), .A1N(n5144), 
        .Y(n2858) );
  OAI2BB2X1 U7271 ( .B0(n5038), .B1(n5529), .A0N(w_matrix[705]), .A1N(n5155), 
        .Y(n2730) );
  OAI2BB2X1 U7272 ( .B0(n5027), .B1(n5407), .A0N(w_matrix[2]), .A1N(n5092), 
        .Y(n3433) );
  OAI2BB2X1 U7273 ( .B0(n5027), .B1(n5429), .A0N(w_matrix[130]), .A1N(n5102), 
        .Y(n3305) );
  OAI2BB2X1 U7274 ( .B0(n5027), .B1(n5506), .A0N(w_matrix[578]), .A1N(n5144), 
        .Y(n2857) );
  OAI2BB2X1 U7275 ( .B0(n5027), .B1(n5529), .A0N(w_matrix[706]), .A1N(n5155), 
        .Y(n2729) );
  OAI2BB2X1 U7276 ( .B0(n5016), .B1(n5407), .A0N(w_matrix[3]), .A1N(n5092), 
        .Y(n3432) );
  OAI2BB2X1 U7277 ( .B0(n5016), .B1(n5429), .A0N(w_matrix[131]), .A1N(n5102), 
        .Y(n3304) );
  OAI2BB2X1 U7278 ( .B0(n5016), .B1(n5506), .A0N(w_matrix[579]), .A1N(n5144), 
        .Y(n2856) );
  OAI2BB2X1 U7279 ( .B0(n5016), .B1(n5529), .A0N(w_matrix[707]), .A1N(n5155), 
        .Y(n2728) );
  OAI2BB2X1 U7280 ( .B0(n5005), .B1(n5407), .A0N(w_matrix[4]), .A1N(n5092), 
        .Y(n3431) );
  OAI2BB2X1 U7281 ( .B0(n5005), .B1(n5429), .A0N(w_matrix[132]), .A1N(n5102), 
        .Y(n3303) );
  OAI2BB2X1 U7282 ( .B0(n5005), .B1(n5506), .A0N(w_matrix[580]), .A1N(n5144), 
        .Y(n2855) );
  OAI2BB2X1 U7283 ( .B0(n5005), .B1(n5529), .A0N(w_matrix[708]), .A1N(n5155), 
        .Y(n2727) );
  OAI2BB2X1 U7284 ( .B0(n4994), .B1(n5407), .A0N(w_matrix[5]), .A1N(n5092), 
        .Y(n3430) );
  OAI2BB2X1 U7285 ( .B0(n4994), .B1(n5429), .A0N(w_matrix[133]), .A1N(n5102), 
        .Y(n3302) );
  OAI2BB2X1 U7286 ( .B0(n4994), .B1(n5506), .A0N(w_matrix[581]), .A1N(n5144), 
        .Y(n2854) );
  OAI2BB2X1 U7287 ( .B0(n4994), .B1(n5529), .A0N(w_matrix[709]), .A1N(n5155), 
        .Y(n2726) );
  OAI2BB2X1 U7288 ( .B0(n4989), .B1(n5407), .A0N(w_matrix[6]), .A1N(n5092), 
        .Y(n3429) );
  OAI2BB2X1 U7289 ( .B0(n4989), .B1(n5429), .A0N(w_matrix[134]), .A1N(n5102), 
        .Y(n3301) );
  OAI2BB2X1 U7290 ( .B0(n4989), .B1(n5506), .A0N(w_matrix[582]), .A1N(n5144), 
        .Y(n2853) );
  OAI2BB2X1 U7291 ( .B0(n4989), .B1(n5529), .A0N(w_matrix[710]), .A1N(n5155), 
        .Y(n2725) );
  OAI2BB2X1 U7292 ( .B0(n4988), .B1(n5407), .A0N(w_matrix[7]), .A1N(n5092), 
        .Y(n3428) );
  OAI2BB2X1 U7293 ( .B0(n4988), .B1(n5429), .A0N(w_matrix[135]), .A1N(n5102), 
        .Y(n3300) );
  OAI2BB2X1 U7294 ( .B0(n4988), .B1(n5506), .A0N(w_matrix[583]), .A1N(n5144), 
        .Y(n2852) );
  OAI2BB2X1 U7295 ( .B0(n4988), .B1(n5529), .A0N(w_matrix[711]), .A1N(n5155), 
        .Y(n2724) );
  OAI2BB2X1 U7296 ( .B0(n4987), .B1(n5407), .A0N(w_matrix[8]), .A1N(n5092), 
        .Y(n3427) );
  OAI2BB2X1 U7297 ( .B0(n4987), .B1(n5429), .A0N(w_matrix[136]), .A1N(n5102), 
        .Y(n3299) );
  OAI2BB2X1 U7298 ( .B0(n4987), .B1(n5506), .A0N(w_matrix[584]), .A1N(n5144), 
        .Y(n2851) );
  OAI2BB2X1 U7299 ( .B0(n4987), .B1(n5529), .A0N(w_matrix[712]), .A1N(n5155), 
        .Y(n2723) );
  OAI2BB2X1 U7300 ( .B0(n4999), .B1(n5416), .A0N(w_matrix[119]), .A1N(n5342), 
        .Y(n3316) );
  OAI2BB2X1 U7301 ( .B0(n4999), .B1(n5438), .A0N(w_matrix[247]), .A1N(n5355), 
        .Y(n3188) );
  OAI2BB2X1 U7302 ( .B0(n4998), .B1(n5416), .A0N(w_matrix[120]), .A1N(n5339), 
        .Y(n3315) );
  OAI2BB2X1 U7303 ( .B0(n4998), .B1(n5438), .A0N(w_matrix[248]), .A1N(n5352), 
        .Y(n3187) );
  OAI2BB2X1 U7304 ( .B0(n4997), .B1(n5416), .A0N(w_matrix[121]), .A1N(n5343), 
        .Y(n3314) );
  OAI2BB2X1 U7305 ( .B0(n4997), .B1(n5438), .A0N(w_matrix[249]), .A1N(n5356), 
        .Y(n3186) );
  OAI2BB2X1 U7306 ( .B0(n4996), .B1(n5416), .A0N(w_matrix[122]), .A1N(n5344), 
        .Y(n3313) );
  OAI2BB2X1 U7307 ( .B0(n4996), .B1(n5438), .A0N(w_matrix[250]), .A1N(n5357), 
        .Y(n3185) );
  OAI2BB2X1 U7308 ( .B0(n4995), .B1(n5416), .A0N(w_matrix[123]), .A1N(n5345), 
        .Y(n3312) );
  OAI2BB2X1 U7309 ( .B0(n4995), .B1(n5438), .A0N(w_matrix[251]), .A1N(n5358), 
        .Y(n3184) );
  OAI2BB2X1 U7310 ( .B0(n4993), .B1(n5416), .A0N(w_matrix[124]), .A1N(n5346), 
        .Y(n3311) );
  OAI2BB2X1 U7311 ( .B0(n4993), .B1(n5438), .A0N(w_matrix[252]), .A1N(n5359), 
        .Y(n3183) );
  OAI2BB2X1 U7312 ( .B0(n4992), .B1(n5416), .A0N(w_matrix[125]), .A1N(n5346), 
        .Y(n3310) );
  OAI2BB2X1 U7313 ( .B0(n4992), .B1(n5438), .A0N(w_matrix[253]), .A1N(n5359), 
        .Y(n3182) );
  OAI2BB2X1 U7314 ( .B0(n4991), .B1(n5416), .A0N(w_matrix[126]), .A1N(n5341), 
        .Y(n3309) );
  OAI2BB2X1 U7315 ( .B0(n4991), .B1(n5438), .A0N(w_matrix[254]), .A1N(n5354), 
        .Y(n3181) );
  OAI2BB2X1 U7316 ( .B0(n4990), .B1(n5416), .A0N(w_matrix[127]), .A1N(n5342), 
        .Y(n3308) );
  OAI2BB2X1 U7317 ( .B0(n4990), .B1(n5438), .A0N(w_matrix[255]), .A1N(n5355), 
        .Y(n3180) );
  OAI2BB2X1 U7318 ( .B0(n5045), .B1(n5420), .A0N(w_matrix[77]), .A1N(n5345), 
        .Y(n3358) );
  OAI2BB2X1 U7319 ( .B0(n5045), .B1(n5442), .A0N(w_matrix[205]), .A1N(n5358), 
        .Y(n3230) );
  OAI2BB2X1 U7320 ( .B0(n5044), .B1(n5420), .A0N(w_matrix[78]), .A1N(n5346), 
        .Y(n3357) );
  OAI2BB2X1 U7321 ( .B0(n5044), .B1(n5442), .A0N(w_matrix[206]), .A1N(n5359), 
        .Y(n3229) );
  OAI2BB2X1 U7322 ( .B0(n5043), .B1(n5420), .A0N(w_matrix[79]), .A1N(n5340), 
        .Y(n3356) );
  OAI2BB2X1 U7323 ( .B0(n5043), .B1(n5442), .A0N(w_matrix[207]), .A1N(n5353), 
        .Y(n3228) );
  OAI2BB2X1 U7324 ( .B0(n5001), .B1(n5493), .A0N(w_matrix[565]), .A1N(n5366), 
        .Y(n2870) );
  OAI2BB2X1 U7325 ( .B0(n5001), .B1(n5515), .A0N(w_matrix[693]), .A1N(n5388), 
        .Y(n2742) );
  OAI2BB2X1 U7326 ( .B0(n4999), .B1(n5493), .A0N(w_matrix[567]), .A1N(n5366), 
        .Y(n2868) );
  OAI2BB2X1 U7327 ( .B0(n4999), .B1(n5515), .A0N(w_matrix[695]), .A1N(n5388), 
        .Y(n2740) );
  OAI2BB2X1 U7328 ( .B0(n4997), .B1(n5493), .A0N(w_matrix[569]), .A1N(n5367), 
        .Y(n2866) );
  OAI2BB2X1 U7329 ( .B0(n4997), .B1(n5515), .A0N(w_matrix[697]), .A1N(n5389), 
        .Y(n2738) );
  OAI2BB2X1 U7330 ( .B0(n4995), .B1(n5493), .A0N(w_matrix[571]), .A1N(n5367), 
        .Y(n2864) );
  OAI2BB2X1 U7331 ( .B0(n4995), .B1(n5515), .A0N(w_matrix[699]), .A1N(n5389), 
        .Y(n2736) );
  OAI2BB2X1 U7332 ( .B0(n4992), .B1(n5493), .A0N(w_matrix[573]), .A1N(n5367), 
        .Y(n2862) );
  OAI2BB2X1 U7333 ( .B0(n4992), .B1(n5515), .A0N(w_matrix[701]), .A1N(n5389), 
        .Y(n2734) );
  OAI2BB2X1 U7334 ( .B0(n5049), .B1(n5497), .A0N(w_matrix[512]), .A1N(n5362), 
        .Y(n2923) );
  OAI2BB2X1 U7335 ( .B0(n5049), .B1(n5519), .A0N(w_matrix[640]), .A1N(n5384), 
        .Y(n2795) );
  OAI2BB2X1 U7336 ( .B0(n5038), .B1(n5497), .A0N(w_matrix[513]), .A1N(n5362), 
        .Y(n2922) );
  OAI2BB2X1 U7337 ( .B0(n5038), .B1(n5519), .A0N(w_matrix[641]), .A1N(n5384), 
        .Y(n2794) );
  OAI2BB2X1 U7338 ( .B0(n5027), .B1(n5497), .A0N(w_matrix[514]), .A1N(n5362), 
        .Y(n2921) );
  OAI2BB2X1 U7339 ( .B0(n5027), .B1(n5519), .A0N(w_matrix[642]), .A1N(n5384), 
        .Y(n2793) );
  OAI2BB2X1 U7340 ( .B0(n5016), .B1(n5497), .A0N(w_matrix[515]), .A1N(n5362), 
        .Y(n2920) );
  OAI2BB2X1 U7341 ( .B0(n5016), .B1(n5519), .A0N(w_matrix[643]), .A1N(n5384), 
        .Y(n2792) );
  OAI2BB2X1 U7342 ( .B0(n5005), .B1(n5497), .A0N(w_matrix[516]), .A1N(n5362), 
        .Y(n2919) );
  OAI2BB2X1 U7343 ( .B0(n5005), .B1(n5519), .A0N(w_matrix[644]), .A1N(n5384), 
        .Y(n2791) );
  OAI2BB2X1 U7344 ( .B0(n4994), .B1(n5497), .A0N(w_matrix[517]), .A1N(n5363), 
        .Y(n2918) );
  OAI2BB2X1 U7345 ( .B0(n4994), .B1(n5519), .A0N(w_matrix[645]), .A1N(n5385), 
        .Y(n2790) );
  OAI2BB2X1 U7346 ( .B0(n4989), .B1(n5497), .A0N(w_matrix[518]), .A1N(n5363), 
        .Y(n2917) );
  OAI2BB2X1 U7347 ( .B0(n4989), .B1(n5519), .A0N(w_matrix[646]), .A1N(n5385), 
        .Y(n2789) );
  OAI222XL U7348 ( .A0(n5570), .A1(n4985), .B0(n5565), .B1(n4960), .C0(n5559), 
        .C1(n5929), .Y(n3595) );
  INVX1 U7349 ( .A(x_matrix[624]), .Y(n5929) );
  OAI222XL U7350 ( .A0(n5570), .A1(n4984), .B0(n5566), .B1(n4949), .C0(n5561), 
        .C1(n5928), .Y(n3585) );
  INVX1 U7351 ( .A(x_matrix[634]), .Y(n5928) );
  OAI222XL U7352 ( .A0(n5570), .A1(n4983), .B0(n5565), .B1(n4948), .C0(n5561), 
        .C1(n5927), .Y(n3584) );
  INVX1 U7353 ( .A(x_matrix[635]), .Y(n5927) );
  OAI222XL U7354 ( .A0(n5570), .A1(n4982), .B0(n5564), .B1(n4947), .C0(n5561), 
        .C1(n5926), .Y(n3583) );
  INVX1 U7355 ( .A(x_matrix[636]), .Y(n5926) );
  OAI222XL U7356 ( .A0(n5569), .A1(n4981), .B0(n5564), .B1(n4946), .C0(n5561), 
        .C1(n5925), .Y(n3582) );
  INVX1 U7357 ( .A(x_matrix[637]), .Y(n5925) );
  OAI222XL U7358 ( .A0(n5569), .A1(n4980), .B0(n5564), .B1(n4945), .C0(n5561), 
        .C1(n5924), .Y(n3581) );
  INVX1 U7359 ( .A(x_matrix[638]), .Y(n5924) );
  OAI222XL U7360 ( .A0(n5569), .A1(n4979), .B0(n5564), .B1(n4944), .C0(n5561), 
        .C1(n5923), .Y(n3580) );
  INVX1 U7361 ( .A(x_matrix[639]), .Y(n5923) );
  OAI222XL U7362 ( .A0(n5570), .A1(n4974), .B0(n5566), .B1(n4959), .C0(n5562), 
        .C1(n5918), .Y(n3594) );
  INVX1 U7363 ( .A(x_matrix[625]), .Y(n5918) );
  OAI222XL U7364 ( .A0(n5570), .A1(n4963), .B0(n5565), .B1(n4958), .C0(n5562), 
        .C1(n5907), .Y(n3593) );
  INVX1 U7365 ( .A(x_matrix[626]), .Y(n5907) );
  OAI222XL U7366 ( .A0(n5570), .A1(n4952), .B0(n5566), .B1(n4957), .C0(n5562), 
        .C1(n5904), .Y(n3592) );
  INVX1 U7367 ( .A(x_matrix[627]), .Y(n5904) );
  OAI222XL U7368 ( .A0(n5570), .A1(n4941), .B0(n5564), .B1(n4956), .C0(n5561), 
        .C1(n5903), .Y(n3591) );
  INVX1 U7369 ( .A(x_matrix[628]), .Y(n5903) );
  OAI222XL U7370 ( .A0(n5570), .A1(n4930), .B0(n5565), .B1(n4955), .C0(n5561), 
        .C1(n5902), .Y(n3590) );
  INVX1 U7371 ( .A(x_matrix[629]), .Y(n5902) );
  OAI222XL U7372 ( .A0(n5570), .A1(n4925), .B0(n5566), .B1(n4954), .C0(n5561), 
        .C1(n5901), .Y(n3589) );
  INVX1 U7373 ( .A(x_matrix[630]), .Y(n5901) );
  OAI222XL U7374 ( .A0(n5570), .A1(n4924), .B0(n5564), .B1(n4953), .C0(n5561), 
        .C1(n5900), .Y(n3588) );
  INVX1 U7375 ( .A(x_matrix[631]), .Y(n5900) );
  OAI222XL U7376 ( .A0(n5570), .A1(n4923), .B0(n5565), .B1(n4951), .C0(n5561), 
        .C1(n5899), .Y(n3587) );
  INVX1 U7377 ( .A(x_matrix[632]), .Y(n5899) );
  OAI222XL U7378 ( .A0(n5570), .A1(n4922), .B0(n5564), .B1(n4950), .C0(n5561), 
        .C1(n5898), .Y(n3586) );
  INVX1 U7379 ( .A(x_matrix[633]), .Y(n5898) );
  OAI222XL U7380 ( .A0(n5566), .A1(n4943), .B0(n5569), .B1(n4978), .C0(n5561), 
        .C1(n5922), .Y(n3579) );
  INVX1 U7381 ( .A(x_matrix[640]), .Y(n5922) );
  OAI222XL U7382 ( .A0(n5566), .A1(n4942), .B0(n5569), .B1(n4977), .C0(n5561), 
        .C1(n5921), .Y(n3578) );
  INVX1 U7383 ( .A(x_matrix[641]), .Y(n5921) );
  OAI222XL U7384 ( .A0(n5566), .A1(n4940), .B0(n5569), .B1(n4976), .C0(n5562), 
        .C1(n5920), .Y(n3577) );
  INVX1 U7385 ( .A(x_matrix[642]), .Y(n5920) );
  OAI222XL U7386 ( .A0(n5566), .A1(n4939), .B0(n5569), .B1(n4975), .C0(n5561), 
        .C1(n5919), .Y(n3576) );
  INVX1 U7387 ( .A(x_matrix[643]), .Y(n5919) );
  OAI222XL U7388 ( .A0(n5566), .A1(n4938), .B0(n5569), .B1(n4973), .C0(n5560), 
        .C1(n5917), .Y(n3575) );
  INVX1 U7389 ( .A(x_matrix[644]), .Y(n5917) );
  OAI222XL U7390 ( .A0(n5566), .A1(n4937), .B0(n5569), .B1(n4972), .C0(n5560), 
        .C1(n5916), .Y(n3574) );
  INVX1 U7391 ( .A(x_matrix[645]), .Y(n5916) );
  OAI222XL U7392 ( .A0(n5566), .A1(n4936), .B0(n5569), .B1(n4971), .C0(n5560), 
        .C1(n5915), .Y(n3573) );
  INVX1 U7393 ( .A(x_matrix[646]), .Y(n5915) );
  OAI222XL U7394 ( .A0(n5566), .A1(n4935), .B0(n5569), .B1(n4970), .C0(n5560), 
        .C1(n5914), .Y(n3572) );
  INVX1 U7395 ( .A(x_matrix[647]), .Y(n5914) );
  OAI222XL U7396 ( .A0(n5566), .A1(n4934), .B0(n5569), .B1(n4969), .C0(n5560), 
        .C1(n5913), .Y(n3571) );
  INVX1 U7397 ( .A(x_matrix[648]), .Y(n5913) );
  OAI222XL U7398 ( .A0(n5566), .A1(n4933), .B0(n5569), .B1(n4968), .C0(n5560), 
        .C1(n5912), .Y(n3570) );
  INVX1 U7399 ( .A(x_matrix[649]), .Y(n5912) );
  OAI222XL U7400 ( .A0(n5566), .A1(n4932), .B0(n5569), .B1(n4967), .C0(n5562), 
        .C1(n5911), .Y(n3569) );
  INVX1 U7401 ( .A(x_matrix[650]), .Y(n5911) );
  OAI222XL U7402 ( .A0(n5566), .A1(n4931), .B0(n5569), .B1(n4966), .C0(n5560), 
        .C1(n5910), .Y(n3568) );
  INVX1 U7403 ( .A(x_matrix[651]), .Y(n5910) );
  OAI222XL U7404 ( .A0(n5566), .A1(n4929), .B0(n5569), .B1(n4965), .C0(n5560), 
        .C1(n5909), .Y(n3567) );
  INVX1 U7405 ( .A(x_matrix[652]), .Y(n5909) );
  OAI222XL U7406 ( .A0(n5565), .A1(n4928), .B0(n5569), .B1(n4964), .C0(n5562), 
        .C1(n5908), .Y(n3566) );
  INVX1 U7407 ( .A(x_matrix[653]), .Y(n5908) );
  OAI222XL U7408 ( .A0(n5565), .A1(n4927), .B0(n5569), .B1(n4962), .C0(n5560), 
        .C1(n5906), .Y(n3565) );
  INVX1 U7409 ( .A(x_matrix[654]), .Y(n5906) );
  OAI222XL U7410 ( .A0(n5565), .A1(n4926), .B0(n5569), .B1(n4961), .C0(n5562), 
        .C1(n5905), .Y(n3564) );
  INVX1 U7411 ( .A(x_matrix[655]), .Y(n5905) );
  OAI222XL U7412 ( .A0(n5049), .A1(n5569), .B0(n5024), .B1(n5564), .C0(n5559), 
        .C1(n673), .Y(n2571) );
  OAI222X1 U7413 ( .A0(n5048), .A1(n5569), .B0(n5013), .B1(n5564), .C0(n5560), 
        .C1(n663), .Y(n2561) );
  OAI222X1 U7414 ( .A0(n5047), .A1(n5569), .B0(n5012), .B1(n5566), .C0(n5559), 
        .C1(n662), .Y(n2560) );
  OAI222X1 U7415 ( .A0(n5046), .A1(n5569), .B0(n5011), .B1(n5565), .C0(n5559), 
        .C1(n661), .Y(n2559) );
  OAI222X1 U7416 ( .A0(n5045), .A1(n5569), .B0(n5010), .B1(n5566), .C0(n5559), 
        .C1(n660), .Y(n2558) );
  OAI222X1 U7417 ( .A0(n5044), .A1(n5569), .B0(n5009), .B1(n5564), .C0(n5559), 
        .C1(n659), .Y(n2557) );
  OAI222X1 U7418 ( .A0(n5043), .A1(n5569), .B0(n5008), .B1(n5564), .C0(n5560), 
        .C1(n658), .Y(n2556) );
  OAI222X1 U7419 ( .A0(n5038), .A1(n5569), .B0(n5023), .B1(n5564), .C0(n5561), 
        .C1(n672), .Y(n2570) );
  OAI222X1 U7420 ( .A0(n5027), .A1(n5569), .B0(n5022), .B1(n5564), .C0(n5561), 
        .C1(n671), .Y(n2569) );
  OAI222X1 U7421 ( .A0(n5016), .A1(n5569), .B0(n5021), .B1(n5564), .C0(n5560), 
        .C1(n670), .Y(n2568) );
  OAI222X1 U7422 ( .A0(n5005), .A1(n5569), .B0(n5020), .B1(n889), .C0(n5560), 
        .C1(n669), .Y(n2567) );
  OAI222X1 U7423 ( .A0(n4994), .A1(n5569), .B0(n5019), .B1(n5564), .C0(n5560), 
        .C1(n668), .Y(n2566) );
  OAI222X1 U7424 ( .A0(n4989), .A1(n5569), .B0(n5018), .B1(n5564), .C0(n5560), 
        .C1(n667), .Y(n2565) );
  OAI222X1 U7425 ( .A0(n4988), .A1(n5569), .B0(n5017), .B1(n889), .C0(n5560), 
        .C1(n666), .Y(n2564) );
  OAI222X1 U7426 ( .A0(n4987), .A1(n5569), .B0(n5015), .B1(n889), .C0(n5560), 
        .C1(n665), .Y(n2563) );
  OAI222X1 U7427 ( .A0(n4986), .A1(n5569), .B0(n5014), .B1(n889), .C0(n5560), 
        .C1(n664), .Y(n2562) );
  OAI221XL U7428 ( .A0(n5042), .A1(n5569), .B0(n5007), .B1(n5565), .C0(n905), 
        .Y(n2555) );
  NAND2X1 U7429 ( .A(w_matrix[880]), .B(n5558), .Y(n905) );
  OAI221XL U7430 ( .A0(n5041), .A1(n5569), .B0(n5006), .B1(n5565), .C0(n904), 
        .Y(n2554) );
  NAND2X1 U7431 ( .A(w_matrix[881]), .B(n5558), .Y(n904) );
  OAI221XL U7432 ( .A0(n5040), .A1(n5569), .B0(n5004), .B1(n5565), .C0(n903), 
        .Y(n2553) );
  NAND2X1 U7433 ( .A(w_matrix[882]), .B(n5558), .Y(n903) );
  OAI221XL U7434 ( .A0(n5039), .A1(n5569), .B0(n5003), .B1(n5565), .C0(n902), 
        .Y(n2552) );
  NAND2X1 U7435 ( .A(w_matrix[883]), .B(n5558), .Y(n902) );
  OAI221XL U7436 ( .A0(n5037), .A1(n5569), .B0(n5002), .B1(n5565), .C0(n901), 
        .Y(n2551) );
  NAND2X1 U7437 ( .A(w_matrix[884]), .B(n5558), .Y(n901) );
  OAI221XL U7438 ( .A0(n5036), .A1(n5569), .B0(n5001), .B1(n5565), .C0(n900), 
        .Y(n2550) );
  NAND2X1 U7439 ( .A(w_matrix[885]), .B(n5558), .Y(n900) );
  OAI221XL U7440 ( .A0(n5035), .A1(n5569), .B0(n5000), .B1(n5564), .C0(n899), 
        .Y(n2549) );
  NAND2X1 U7441 ( .A(w_matrix[886]), .B(n5558), .Y(n899) );
  OAI221XL U7442 ( .A0(n5034), .A1(n5569), .B0(n4999), .B1(n5564), .C0(n898), 
        .Y(n2548) );
  NAND2X1 U7443 ( .A(w_matrix[887]), .B(n5558), .Y(n898) );
  OAI221XL U7444 ( .A0(n5033), .A1(n5569), .B0(n4998), .B1(n5565), .C0(n897), 
        .Y(n2547) );
  NAND2X1 U7445 ( .A(w_matrix[888]), .B(n5558), .Y(n897) );
  OAI221XL U7446 ( .A0(n5032), .A1(n5569), .B0(n4997), .B1(n5564), .C0(n896), 
        .Y(n2546) );
  NAND2X1 U7447 ( .A(w_matrix[889]), .B(n5558), .Y(n896) );
  OAI221XL U7448 ( .A0(n5031), .A1(n5569), .B0(n4996), .B1(n5564), .C0(n895), 
        .Y(n2545) );
  NAND2X1 U7449 ( .A(w_matrix[890]), .B(n5558), .Y(n895) );
  OAI221XL U7450 ( .A0(n5030), .A1(n5569), .B0(n4995), .B1(n5565), .C0(n894), 
        .Y(n2544) );
  NAND2X1 U7451 ( .A(w_matrix[891]), .B(n5558), .Y(n894) );
  OAI221XL U7452 ( .A0(n5029), .A1(n5569), .B0(n4993), .B1(n5565), .C0(n893), 
        .Y(n2543) );
  NAND2X1 U7453 ( .A(w_matrix[892]), .B(n5558), .Y(n893) );
  OAI221XL U7454 ( .A0(n5028), .A1(n5569), .B0(n4992), .B1(n5566), .C0(n892), 
        .Y(n2542) );
  NAND2X1 U7455 ( .A(w_matrix[893]), .B(n5558), .Y(n892) );
  OAI221XL U7456 ( .A0(n5026), .A1(n5569), .B0(n4991), .B1(n5565), .C0(n891), 
        .Y(n2541) );
  NAND2X1 U7457 ( .A(w_matrix[894]), .B(n5558), .Y(n891) );
  OAI221XL U7458 ( .A0(n5025), .A1(n5569), .B0(n4990), .B1(n5565), .C0(n890), 
        .Y(n2540) );
  NAND2X1 U7459 ( .A(w_matrix[895]), .B(n5558), .Y(n890) );
  OAI2BB2X1 U7460 ( .B0(n5049), .B1(n5554), .A0N(w_matrix[832]), .A1N(n5548), 
        .Y(n2603) );
  OAI2BB2X1 U7461 ( .B0(n5585), .B1(n5029), .A0N(w_matrix[988]), .A1N(n5181), 
        .Y(n2447) );
  OAI2BB2X1 U7462 ( .B0(n5585), .B1(n5028), .A0N(w_matrix[989]), .A1N(n5181), 
        .Y(n2446) );
  OAI2BB2X1 U7463 ( .B0(n5583), .B1(n5026), .A0N(w_matrix[990]), .A1N(n5181), 
        .Y(n2445) );
  OAI2BB2X1 U7464 ( .B0(n5584), .B1(n5025), .A0N(w_matrix[991]), .A1N(n5178), 
        .Y(n2444) );
  OAI2BB2X1 U7465 ( .B0(n5591), .B1(n4993), .A0N(w_matrix[1020]), .A1N(n5187), 
        .Y(n2415) );
  OAI2BB2X1 U7466 ( .B0(n5591), .B1(n4992), .A0N(w_matrix[1021]), .A1N(n5187), 
        .Y(n2414) );
  OAI2BB2X1 U7467 ( .B0(n5589), .B1(n4991), .A0N(w_matrix[1022]), .A1N(n5187), 
        .Y(n2413) );
  OAI2BB2X1 U7468 ( .B0(n5590), .B1(n4990), .A0N(w_matrix[1023]), .A1N(n5183), 
        .Y(n2412) );
  OAI2BB2X1 U7469 ( .B0(n5552), .B1(n4985), .A0N(n5547), .A1N(x_matrix[592]), 
        .Y(n3627) );
  OAI2BB2X1 U7470 ( .B0(n5582), .B1(n4985), .A0N(n5177), .A1N(x_matrix[704]), 
        .Y(n3499) );
  OAI2BB2X1 U7471 ( .B0(n5552), .B1(n4984), .A0N(n5547), .A1N(x_matrix[602]), 
        .Y(n3617) );
  OAI2BB2X1 U7472 ( .B0(n5582), .B1(n4984), .A0N(n5177), .A1N(x_matrix[714]), 
        .Y(n3489) );
  OAI2BB2X1 U7473 ( .B0(n5552), .B1(n4983), .A0N(n5548), .A1N(x_matrix[603]), 
        .Y(n3616) );
  OAI2BB2X1 U7474 ( .B0(n5582), .B1(n4983), .A0N(n5177), .A1N(x_matrix[715]), 
        .Y(n3488) );
  OAI2BB2X1 U7475 ( .B0(n5552), .B1(n4982), .A0N(n5547), .A1N(x_matrix[604]), 
        .Y(n3615) );
  OAI2BB2X1 U7476 ( .B0(n5582), .B1(n4982), .A0N(n5178), .A1N(x_matrix[716]), 
        .Y(n3487) );
  OAI2BB2X1 U7477 ( .B0(n5552), .B1(n4981), .A0N(n5547), .A1N(x_matrix[605]), 
        .Y(n3614) );
  OAI2BB2X1 U7478 ( .B0(n5585), .B1(n4981), .A0N(n5178), .A1N(x_matrix[717]), 
        .Y(n3486) );
  OAI2BB2X1 U7479 ( .B0(n5552), .B1(n4980), .A0N(n5547), .A1N(x_matrix[606]), 
        .Y(n3613) );
  OAI2BB2X1 U7480 ( .B0(n5582), .B1(n4980), .A0N(n5178), .A1N(x_matrix[718]), 
        .Y(n3485) );
  OAI2BB2X1 U7481 ( .B0(n5552), .B1(n4979), .A0N(n5547), .A1N(x_matrix[607]), 
        .Y(n3612) );
  OAI2BB2X1 U7482 ( .B0(n5582), .B1(n4979), .A0N(n5178), .A1N(x_matrix[719]), 
        .Y(n3484) );
  OAI2BB2X1 U7483 ( .B0(n5552), .B1(n4974), .A0N(n908), .A1N(x_matrix[593]), 
        .Y(n3626) );
  OAI2BB2X1 U7484 ( .B0(n5582), .B1(n4974), .A0N(n5177), .A1N(x_matrix[705]), 
        .Y(n3498) );
  OAI2BB2X1 U7485 ( .B0(n5552), .B1(n4963), .A0N(n908), .A1N(x_matrix[594]), 
        .Y(n3625) );
  OAI2BB2X1 U7486 ( .B0(n5582), .B1(n4963), .A0N(n5177), .A1N(x_matrix[706]), 
        .Y(n3497) );
  OAI2BB2X1 U7487 ( .B0(n5552), .B1(n4952), .A0N(n908), .A1N(x_matrix[595]), 
        .Y(n3624) );
  OAI2BB2X1 U7488 ( .B0(n5582), .B1(n4952), .A0N(n5177), .A1N(x_matrix[707]), 
        .Y(n3496) );
  OAI2BB2X1 U7489 ( .B0(n5552), .B1(n4941), .A0N(n908), .A1N(x_matrix[596]), 
        .Y(n3623) );
  OAI2BB2X1 U7490 ( .B0(n5582), .B1(n4941), .A0N(n5177), .A1N(x_matrix[708]), 
        .Y(n3495) );
  OAI2BB2X1 U7491 ( .B0(n5552), .B1(n4930), .A0N(n908), .A1N(x_matrix[597]), 
        .Y(n3622) );
  OAI2BB2X1 U7492 ( .B0(n5582), .B1(n4930), .A0N(n5177), .A1N(x_matrix[709]), 
        .Y(n3494) );
  OAI2BB2X1 U7493 ( .B0(n5552), .B1(n4925), .A0N(n908), .A1N(x_matrix[598]), 
        .Y(n3621) );
  OAI2BB2X1 U7494 ( .B0(n5582), .B1(n4925), .A0N(n5177), .A1N(x_matrix[710]), 
        .Y(n3493) );
  OAI2BB2X1 U7495 ( .B0(n5552), .B1(n4924), .A0N(n908), .A1N(x_matrix[599]), 
        .Y(n3620) );
  OAI2BB2X1 U7496 ( .B0(n5582), .B1(n4924), .A0N(n5177), .A1N(x_matrix[711]), 
        .Y(n3492) );
  OAI2BB2X1 U7497 ( .B0(n5552), .B1(n4923), .A0N(n908), .A1N(x_matrix[600]), 
        .Y(n3619) );
  OAI2BB2X1 U7498 ( .B0(n5582), .B1(n4923), .A0N(n5177), .A1N(x_matrix[712]), 
        .Y(n3491) );
  OAI2BB2X1 U7499 ( .B0(n5552), .B1(n4922), .A0N(n908), .A1N(x_matrix[601]), 
        .Y(n3618) );
  OAI2BB2X1 U7500 ( .B0(n5582), .B1(n4922), .A0N(n5177), .A1N(x_matrix[713]), 
        .Y(n3490) );
  OAI2BB2X1 U7501 ( .B0(n5553), .B1(n4978), .A0N(n5547), .A1N(x_matrix[608]), 
        .Y(n3611) );
  OAI2BB2X1 U7502 ( .B0(n5582), .B1(n4978), .A0N(n5178), .A1N(x_matrix[720]), 
        .Y(n3483) );
  OAI2BB2X1 U7503 ( .B0(n5552), .B1(n4977), .A0N(n5547), .A1N(x_matrix[609]), 
        .Y(n3610) );
  OAI2BB2X1 U7504 ( .B0(n5583), .B1(n4977), .A0N(n5178), .A1N(x_matrix[721]), 
        .Y(n3482) );
  OAI2BB2X1 U7505 ( .B0(n5553), .B1(n4976), .A0N(n5547), .A1N(x_matrix[610]), 
        .Y(n3609) );
  OAI2BB2X1 U7506 ( .B0(n5582), .B1(n4976), .A0N(n5178), .A1N(x_matrix[722]), 
        .Y(n3481) );
  OAI2BB2X1 U7507 ( .B0(n5554), .B1(n4975), .A0N(n5547), .A1N(x_matrix[611]), 
        .Y(n3608) );
  OAI2BB2X1 U7508 ( .B0(n5583), .B1(n4975), .A0N(n5178), .A1N(x_matrix[723]), 
        .Y(n3480) );
  OAI2BB2X1 U7509 ( .B0(n5555), .B1(n4973), .A0N(n5547), .A1N(x_matrix[612]), 
        .Y(n3607) );
  OAI2BB2X1 U7510 ( .B0(n5584), .B1(n4973), .A0N(n5178), .A1N(x_matrix[724]), 
        .Y(n3479) );
  OAI2BB2X1 U7511 ( .B0(n5553), .B1(n4972), .A0N(n5547), .A1N(x_matrix[613]), 
        .Y(n3606) );
  OAI2BB2X1 U7512 ( .B0(n5585), .B1(n4972), .A0N(n5178), .A1N(x_matrix[725]), 
        .Y(n3478) );
  OAI2BB2X1 U7513 ( .B0(n5554), .B1(n4971), .A0N(n5547), .A1N(x_matrix[614]), 
        .Y(n3605) );
  OAI2BB2X1 U7514 ( .B0(n5583), .B1(n4971), .A0N(n5178), .A1N(x_matrix[726]), 
        .Y(n3477) );
  OAI2BB2X1 U7515 ( .B0(n5555), .B1(n4970), .A0N(n5547), .A1N(x_matrix[615]), 
        .Y(n3604) );
  OAI2BB2X1 U7516 ( .B0(n5584), .B1(n4970), .A0N(n5178), .A1N(x_matrix[727]), 
        .Y(n3476) );
  OAI2BB2X1 U7517 ( .B0(n5553), .B1(n4969), .A0N(n5548), .A1N(x_matrix[616]), 
        .Y(n3603) );
  OAI2BB2X1 U7518 ( .B0(n5583), .B1(n4969), .A0N(n5179), .A1N(x_matrix[728]), 
        .Y(n3475) );
  OAI2BB2X1 U7519 ( .B0(n5553), .B1(n4968), .A0N(n5548), .A1N(x_matrix[617]), 
        .Y(n3602) );
  OAI2BB2X1 U7520 ( .B0(n5583), .B1(n4968), .A0N(n5179), .A1N(x_matrix[729]), 
        .Y(n3474) );
  OAI2BB2X1 U7521 ( .B0(n5553), .B1(n4967), .A0N(n5548), .A1N(x_matrix[618]), 
        .Y(n3601) );
  OAI2BB2X1 U7522 ( .B0(n5583), .B1(n4967), .A0N(n5179), .A1N(x_matrix[730]), 
        .Y(n3473) );
  OAI2BB2X1 U7523 ( .B0(n5553), .B1(n4966), .A0N(n5548), .A1N(x_matrix[619]), 
        .Y(n3600) );
  OAI2BB2X1 U7524 ( .B0(n5583), .B1(n4966), .A0N(n5179), .A1N(x_matrix[731]), 
        .Y(n3472) );
  OAI2BB2X1 U7525 ( .B0(n5553), .B1(n4965), .A0N(n5548), .A1N(x_matrix[620]), 
        .Y(n3599) );
  OAI2BB2X1 U7526 ( .B0(n5583), .B1(n4965), .A0N(n5179), .A1N(x_matrix[732]), 
        .Y(n3471) );
  OAI2BB2X1 U7527 ( .B0(n5553), .B1(n4964), .A0N(n5548), .A1N(x_matrix[621]), 
        .Y(n3598) );
  OAI2BB2X1 U7528 ( .B0(n5583), .B1(n4964), .A0N(n5179), .A1N(x_matrix[733]), 
        .Y(n3470) );
  OAI2BB2X1 U7529 ( .B0(n5553), .B1(n4962), .A0N(n5548), .A1N(x_matrix[622]), 
        .Y(n3597) );
  OAI2BB2X1 U7530 ( .B0(n5583), .B1(n4962), .A0N(n5179), .A1N(x_matrix[734]), 
        .Y(n3469) );
  OAI2BB2X1 U7531 ( .B0(n5553), .B1(n4961), .A0N(n5548), .A1N(x_matrix[623]), 
        .Y(n3596) );
  OAI2BB2X1 U7532 ( .B0(n5583), .B1(n4961), .A0N(n5179), .A1N(x_matrix[735]), 
        .Y(n3468) );
  OAI2BB2X1 U7533 ( .B0(n5585), .B1(n5042), .A0N(w_matrix[976]), .A1N(n5180), 
        .Y(n2459) );
  OAI2BB2X1 U7534 ( .B0(n5585), .B1(n5041), .A0N(w_matrix[977]), .A1N(n5180), 
        .Y(n2458) );
  OAI2BB2X1 U7535 ( .B0(n5585), .B1(n5040), .A0N(w_matrix[978]), .A1N(n5181), 
        .Y(n2457) );
  OAI2BB2X1 U7536 ( .B0(n5585), .B1(n5039), .A0N(w_matrix[979]), .A1N(n5181), 
        .Y(n2456) );
  OAI2BB2X1 U7537 ( .B0(n5585), .B1(n5037), .A0N(w_matrix[980]), .A1N(n5181), 
        .Y(n2455) );
  OAI2BB2X1 U7538 ( .B0(n5585), .B1(n5036), .A0N(w_matrix[981]), .A1N(n5181), 
        .Y(n2454) );
  OAI2BB2X1 U7539 ( .B0(n5585), .B1(n5035), .A0N(w_matrix[982]), .A1N(n5181), 
        .Y(n2453) );
  OAI2BB2X1 U7540 ( .B0(n5585), .B1(n5034), .A0N(w_matrix[983]), .A1N(n5181), 
        .Y(n2452) );
  OAI2BB2X1 U7541 ( .B0(n5585), .B1(n5033), .A0N(w_matrix[984]), .A1N(n5181), 
        .Y(n2451) );
  OAI2BB2X1 U7542 ( .B0(n5585), .B1(n5032), .A0N(w_matrix[985]), .A1N(n5181), 
        .Y(n2450) );
  OAI2BB2X1 U7543 ( .B0(n5585), .B1(n5031), .A0N(w_matrix[986]), .A1N(n5181), 
        .Y(n2449) );
  OAI2BB2X1 U7544 ( .B0(n5585), .B1(n5030), .A0N(w_matrix[987]), .A1N(n5181), 
        .Y(n2448) );
  OAI2BB2X1 U7545 ( .B0(n5583), .B1(n5049), .A0N(w_matrix[960]), .A1N(n5179), 
        .Y(n2475) );
  OAI2BB2X1 U7546 ( .B0(n5584), .B1(n5048), .A0N(w_matrix[970]), .A1N(n5180), 
        .Y(n2465) );
  OAI2BB2X1 U7547 ( .B0(n5584), .B1(n5047), .A0N(w_matrix[971]), .A1N(n5180), 
        .Y(n2464) );
  OAI2BB2X1 U7548 ( .B0(n5584), .B1(n5046), .A0N(w_matrix[972]), .A1N(n5180), 
        .Y(n2463) );
  OAI2BB2X1 U7549 ( .B0(n5584), .B1(n5045), .A0N(w_matrix[973]), .A1N(n5180), 
        .Y(n2462) );
  OAI2BB2X1 U7550 ( .B0(n5584), .B1(n5044), .A0N(w_matrix[974]), .A1N(n5180), 
        .Y(n2461) );
  OAI2BB2X1 U7551 ( .B0(n5584), .B1(n5043), .A0N(w_matrix[975]), .A1N(n5180), 
        .Y(n2460) );
  OAI2BB2X1 U7552 ( .B0(n5583), .B1(n5038), .A0N(w_matrix[961]), .A1N(n5179), 
        .Y(n2474) );
  OAI2BB2X1 U7553 ( .B0(n5583), .B1(n5027), .A0N(w_matrix[962]), .A1N(n5179), 
        .Y(n2473) );
  OAI2BB2X1 U7554 ( .B0(n5583), .B1(n5016), .A0N(w_matrix[963]), .A1N(n5179), 
        .Y(n2472) );
  OAI2BB2X1 U7555 ( .B0(n5584), .B1(n5005), .A0N(w_matrix[964]), .A1N(n5179), 
        .Y(n2471) );
  OAI2BB2X1 U7556 ( .B0(n5584), .B1(n4994), .A0N(w_matrix[965]), .A1N(n5180), 
        .Y(n2470) );
  OAI2BB2X1 U7557 ( .B0(n5584), .B1(n4989), .A0N(w_matrix[966]), .A1N(n5180), 
        .Y(n2469) );
  OAI2BB2X1 U7558 ( .B0(n5584), .B1(n4988), .A0N(w_matrix[967]), .A1N(n5180), 
        .Y(n2468) );
  OAI2BB2X1 U7559 ( .B0(n5584), .B1(n4987), .A0N(w_matrix[968]), .A1N(n5180), 
        .Y(n2467) );
  OAI2BB2X1 U7560 ( .B0(n5584), .B1(n4986), .A0N(w_matrix[969]), .A1N(n5180), 
        .Y(n2466) );
  OAI2BB2X1 U7561 ( .B0(n5588), .B1(n4943), .A0N(n5184), .A1N(x_matrix[752]), 
        .Y(n3451) );
  OAI2BB2X1 U7562 ( .B0(n5591), .B1(n4942), .A0N(n5184), .A1N(x_matrix[753]), 
        .Y(n3450) );
  OAI2BB2X1 U7563 ( .B0(n5588), .B1(n4940), .A0N(n5184), .A1N(x_matrix[754]), 
        .Y(n3449) );
  OAI2BB2X1 U7564 ( .B0(n5588), .B1(n4939), .A0N(n5184), .A1N(x_matrix[755]), 
        .Y(n3448) );
  OAI2BB2X1 U7565 ( .B0(n5588), .B1(n4938), .A0N(n5184), .A1N(x_matrix[756]), 
        .Y(n3447) );
  OAI2BB2X1 U7566 ( .B0(n5589), .B1(n4937), .A0N(n5184), .A1N(x_matrix[757]), 
        .Y(n3446) );
  OAI2BB2X1 U7567 ( .B0(n5588), .B1(n4936), .A0N(n5184), .A1N(x_matrix[758]), 
        .Y(n3445) );
  OAI2BB2X1 U7568 ( .B0(n5589), .B1(n4935), .A0N(n5184), .A1N(x_matrix[759]), 
        .Y(n3444) );
  OAI2BB2X1 U7569 ( .B0(n5589), .B1(n4934), .A0N(n5185), .A1N(x_matrix[760]), 
        .Y(n3443) );
  OAI2BB2X1 U7570 ( .B0(n5589), .B1(n4933), .A0N(n5185), .A1N(x_matrix[761]), 
        .Y(n3442) );
  OAI2BB2X1 U7571 ( .B0(n5589), .B1(n4932), .A0N(n5185), .A1N(x_matrix[762]), 
        .Y(n3441) );
  OAI2BB2X1 U7572 ( .B0(n5589), .B1(n4931), .A0N(n5185), .A1N(x_matrix[763]), 
        .Y(n3440) );
  OAI2BB2X1 U7573 ( .B0(n5589), .B1(n4929), .A0N(n5185), .A1N(x_matrix[764]), 
        .Y(n3439) );
  OAI2BB2X1 U7574 ( .B0(n5589), .B1(n4928), .A0N(n5185), .A1N(x_matrix[765]), 
        .Y(n3438) );
  OAI2BB2X1 U7575 ( .B0(n5589), .B1(n4927), .A0N(n5185), .A1N(x_matrix[766]), 
        .Y(n3437) );
  OAI2BB2X1 U7576 ( .B0(n5589), .B1(n4926), .A0N(n5185), .A1N(x_matrix[767]), 
        .Y(n3436) );
  OAI2BB2X1 U7577 ( .B0(n5588), .B1(n4960), .A0N(n5183), .A1N(x_matrix[736]), 
        .Y(n3467) );
  OAI2BB2X1 U7578 ( .B0(n5588), .B1(n4959), .A0N(n5183), .A1N(x_matrix[737]), 
        .Y(n3466) );
  OAI2BB2X1 U7579 ( .B0(n5588), .B1(n4958), .A0N(n5183), .A1N(x_matrix[738]), 
        .Y(n3465) );
  OAI2BB2X1 U7580 ( .B0(n5588), .B1(n4957), .A0N(n5183), .A1N(x_matrix[739]), 
        .Y(n3464) );
  OAI2BB2X1 U7581 ( .B0(n5588), .B1(n4956), .A0N(n5183), .A1N(x_matrix[740]), 
        .Y(n3463) );
  OAI2BB2X1 U7582 ( .B0(n5588), .B1(n4955), .A0N(n5183), .A1N(x_matrix[741]), 
        .Y(n3462) );
  OAI2BB2X1 U7583 ( .B0(n5588), .B1(n4954), .A0N(n5183), .A1N(x_matrix[742]), 
        .Y(n3461) );
  OAI2BB2X1 U7584 ( .B0(n5588), .B1(n4953), .A0N(n5183), .A1N(x_matrix[743]), 
        .Y(n3460) );
  OAI2BB2X1 U7585 ( .B0(n5588), .B1(n4951), .A0N(n5183), .A1N(x_matrix[744]), 
        .Y(n3459) );
  OAI2BB2X1 U7586 ( .B0(n5588), .B1(n4950), .A0N(n5183), .A1N(x_matrix[745]), 
        .Y(n3458) );
  OAI2BB2X1 U7587 ( .B0(n5588), .B1(n4949), .A0N(n5183), .A1N(x_matrix[746]), 
        .Y(n3457) );
  OAI2BB2X1 U7588 ( .B0(n5588), .B1(n4948), .A0N(n5183), .A1N(x_matrix[747]), 
        .Y(n3456) );
  OAI2BB2X1 U7589 ( .B0(n5590), .B1(n4947), .A0N(n5184), .A1N(x_matrix[748]), 
        .Y(n3455) );
  OAI2BB2X1 U7590 ( .B0(n5591), .B1(n4946), .A0N(n5184), .A1N(x_matrix[749]), 
        .Y(n3454) );
  OAI2BB2X1 U7591 ( .B0(n5589), .B1(n4945), .A0N(n5184), .A1N(x_matrix[750]), 
        .Y(n3453) );
  OAI2BB2X1 U7592 ( .B0(n5590), .B1(n4944), .A0N(n5184), .A1N(x_matrix[751]), 
        .Y(n3452) );
  OAI2BB2X1 U7593 ( .B0(n5589), .B1(n5024), .A0N(w_matrix[992]), .A1N(n5185), 
        .Y(n2443) );
  OAI2BB2X1 U7594 ( .B0(n5589), .B1(n5023), .A0N(w_matrix[993]), .A1N(n5185), 
        .Y(n2442) );
  OAI2BB2X1 U7595 ( .B0(n5589), .B1(n5022), .A0N(w_matrix[994]), .A1N(n5185), 
        .Y(n2441) );
  OAI2BB2X1 U7596 ( .B0(n5589), .B1(n5021), .A0N(w_matrix[995]), .A1N(n5185), 
        .Y(n2440) );
  OAI2BB2X1 U7597 ( .B0(n5590), .B1(n5020), .A0N(w_matrix[996]), .A1N(n5185), 
        .Y(n2439) );
  OAI2BB2X1 U7598 ( .B0(n5590), .B1(n5019), .A0N(w_matrix[997]), .A1N(n5186), 
        .Y(n2438) );
  OAI2BB2X1 U7599 ( .B0(n5590), .B1(n5018), .A0N(w_matrix[998]), .A1N(n5186), 
        .Y(n2437) );
  OAI2BB2X1 U7600 ( .B0(n5590), .B1(n5017), .A0N(w_matrix[999]), .A1N(n5186), 
        .Y(n2436) );
  OAI2BB2X1 U7601 ( .B0(n5590), .B1(n5015), .A0N(w_matrix[1000]), .A1N(n5186), 
        .Y(n2435) );
  OAI2BB2X1 U7602 ( .B0(n5590), .B1(n5014), .A0N(w_matrix[1001]), .A1N(n5186), 
        .Y(n2434) );
  OAI2BB2X1 U7603 ( .B0(n5590), .B1(n5013), .A0N(w_matrix[1002]), .A1N(n5186), 
        .Y(n2433) );
  OAI2BB2X1 U7604 ( .B0(n5590), .B1(n5012), .A0N(w_matrix[1003]), .A1N(n5186), 
        .Y(n2432) );
  OAI2BB2X1 U7605 ( .B0(n5590), .B1(n5011), .A0N(w_matrix[1004]), .A1N(n5186), 
        .Y(n2431) );
  OAI2BB2X1 U7606 ( .B0(n5590), .B1(n5010), .A0N(w_matrix[1005]), .A1N(n5186), 
        .Y(n2430) );
  OAI2BB2X1 U7607 ( .B0(n5590), .B1(n5009), .A0N(w_matrix[1006]), .A1N(n5186), 
        .Y(n2429) );
  OAI2BB2X1 U7608 ( .B0(n5590), .B1(n5008), .A0N(w_matrix[1007]), .A1N(n5186), 
        .Y(n2428) );
  OAI2BB2X1 U7609 ( .B0(n5591), .B1(n5007), .A0N(w_matrix[1008]), .A1N(n5186), 
        .Y(n2427) );
  OAI2BB2X1 U7610 ( .B0(n5591), .B1(n5006), .A0N(w_matrix[1009]), .A1N(n5186), 
        .Y(n2426) );
  OAI2BB2X1 U7611 ( .B0(n5591), .B1(n5004), .A0N(w_matrix[1010]), .A1N(n5187), 
        .Y(n2425) );
  OAI2BB2X1 U7612 ( .B0(n5591), .B1(n5003), .A0N(w_matrix[1011]), .A1N(n5187), 
        .Y(n2424) );
  OAI2BB2X1 U7613 ( .B0(n5591), .B1(n5002), .A0N(w_matrix[1012]), .A1N(n5187), 
        .Y(n2423) );
  OAI2BB2X1 U7614 ( .B0(n5591), .B1(n5001), .A0N(w_matrix[1013]), .A1N(n5187), 
        .Y(n2422) );
  OAI2BB2X1 U7615 ( .B0(n5591), .B1(n5000), .A0N(w_matrix[1014]), .A1N(n5187), 
        .Y(n2421) );
  OAI2BB2X1 U7616 ( .B0(n5591), .B1(n4999), .A0N(w_matrix[1015]), .A1N(n5187), 
        .Y(n2420) );
  OAI2BB2X1 U7617 ( .B0(n5591), .B1(n4998), .A0N(w_matrix[1016]), .A1N(n5187), 
        .Y(n2419) );
  OAI2BB2X1 U7618 ( .B0(n5591), .B1(n4997), .A0N(w_matrix[1017]), .A1N(n5187), 
        .Y(n2418) );
  OAI2BB2X1 U7619 ( .B0(n5591), .B1(n4996), .A0N(w_matrix[1018]), .A1N(n5187), 
        .Y(n2417) );
  OAI2BB2X1 U7620 ( .B0(n5591), .B1(n4995), .A0N(w_matrix[1019]), .A1N(n5187), 
        .Y(n2416) );
  OAI2BB2X1 U7621 ( .B0(n5048), .B1(n5555), .A0N(w_matrix[842]), .A1N(n5549), 
        .Y(n2593) );
  OAI2BB2X1 U7622 ( .B0(n5047), .B1(n5555), .A0N(w_matrix[843]), .A1N(n5549), 
        .Y(n2592) );
  OAI2BB2X1 U7623 ( .B0(n5046), .B1(n5555), .A0N(w_matrix[844]), .A1N(n5549), 
        .Y(n2591) );
  OAI2BB2X1 U7624 ( .B0(n5045), .B1(n5555), .A0N(w_matrix[845]), .A1N(n5549), 
        .Y(n2590) );
  OAI2BB2X1 U7625 ( .B0(n5044), .B1(n5554), .A0N(w_matrix[846]), .A1N(n5549), 
        .Y(n2589) );
  OAI2BB2X1 U7626 ( .B0(n5043), .B1(n5554), .A0N(w_matrix[847]), .A1N(n5549), 
        .Y(n2588) );
  OAI2BB2X1 U7627 ( .B0(n5042), .B1(n5554), .A0N(w_matrix[848]), .A1N(n5549), 
        .Y(n2587) );
  OAI2BB2X1 U7628 ( .B0(n5041), .B1(n5554), .A0N(w_matrix[849]), .A1N(n5549), 
        .Y(n2586) );
  OAI2BB2X1 U7629 ( .B0(n5040), .B1(n5554), .A0N(w_matrix[850]), .A1N(n5550), 
        .Y(n2585) );
  OAI2BB2X1 U7630 ( .B0(n5039), .B1(n5554), .A0N(w_matrix[851]), .A1N(n5550), 
        .Y(n2584) );
  OAI2BB2X1 U7631 ( .B0(n5038), .B1(n5555), .A0N(w_matrix[833]), .A1N(n5548), 
        .Y(n2602) );
  OAI2BB2X1 U7632 ( .B0(n5037), .B1(n5554), .A0N(w_matrix[852]), .A1N(n5550), 
        .Y(n2583) );
  OAI2BB2X1 U7633 ( .B0(n5036), .B1(n5554), .A0N(w_matrix[853]), .A1N(n5550), 
        .Y(n2582) );
  OAI2BB2X1 U7634 ( .B0(n5035), .B1(n5554), .A0N(w_matrix[854]), .A1N(n5550), 
        .Y(n2581) );
  OAI2BB2X1 U7635 ( .B0(n5034), .B1(n5554), .A0N(w_matrix[855]), .A1N(n5550), 
        .Y(n2580) );
  OAI2BB2X1 U7636 ( .B0(n5033), .B1(n5554), .A0N(w_matrix[856]), .A1N(n5550), 
        .Y(n2579) );
  OAI2BB2X1 U7637 ( .B0(n5032), .B1(n5554), .A0N(w_matrix[857]), .A1N(n5550), 
        .Y(n2578) );
  OAI2BB2X1 U7638 ( .B0(n5027), .B1(n5555), .A0N(w_matrix[834]), .A1N(n5548), 
        .Y(n2601) );
  OAI2BB2X1 U7639 ( .B0(n5025), .B1(n5554), .A0N(w_matrix[863]), .A1N(n5547), 
        .Y(n2572) );
  OAI2BB2X1 U7640 ( .B0(n5016), .B1(n5555), .A0N(w_matrix[835]), .A1N(n5548), 
        .Y(n2600) );
  OAI2BB2X1 U7641 ( .B0(n5005), .B1(n5555), .A0N(w_matrix[836]), .A1N(n5548), 
        .Y(n2599) );
  OAI2BB2X1 U7642 ( .B0(n4994), .B1(n5555), .A0N(w_matrix[837]), .A1N(n5549), 
        .Y(n2598) );
  OAI2BB2X1 U7643 ( .B0(n4989), .B1(n5555), .A0N(w_matrix[838]), .A1N(n5549), 
        .Y(n2597) );
  OAI2BB2X1 U7644 ( .B0(n4988), .B1(n5555), .A0N(w_matrix[839]), .A1N(n5549), 
        .Y(n2596) );
  OAI2BB2X1 U7645 ( .B0(n4987), .B1(n5555), .A0N(w_matrix[840]), .A1N(n5549), 
        .Y(n2595) );
  OAI2BB2X1 U7646 ( .B0(n4986), .B1(n5555), .A0N(w_matrix[841]), .A1N(n5549), 
        .Y(n2594) );
  OAI2BB2X1 U7647 ( .B0(n5031), .B1(n5553), .A0N(w_matrix[858]), .A1N(n5550), 
        .Y(n2577) );
  OAI2BB2X1 U7648 ( .B0(n5030), .B1(n5553), .A0N(w_matrix[859]), .A1N(n5550), 
        .Y(n2576) );
  OAI2BB2X1 U7649 ( .B0(n5029), .B1(n5553), .A0N(w_matrix[860]), .A1N(n5550), 
        .Y(n2575) );
  OAI2BB2X1 U7650 ( .B0(n5028), .B1(n5553), .A0N(w_matrix[861]), .A1N(n5550), 
        .Y(n2574) );
  OAI2BB2X1 U7651 ( .B0(n5026), .B1(n5553), .A0N(w_matrix[862]), .A1N(n5550), 
        .Y(n2573) );
  INVX1 U7652 ( .A(n1113), .Y(n5803) );
  AOI22X1 U7653 ( .A0(N1302), .A1(n4474), .B0(in_start_addr[0]), .B1(n5069), 
        .Y(n1113) );
  INVX1 U7654 ( .A(n1104), .Y(n5812) );
  AOI22X1 U7655 ( .A0(N1330), .A1(n5067), .B0(weight_start_addr[0]), .B1(n5069), .Y(n1104) );
  OAI2BB1X1 U7656 ( .A0N(N12245), .A1N(n5062), .B0(n1137), .Y(N12605) );
  AOI22X1 U7657 ( .A0(N12125), .A1(n5327), .B0(N12525), .B1(n5325), .Y(n1137)
         );
  INVX1 U7658 ( .A(n959), .Y(n5796) );
  AOI22X1 U7659 ( .A0(N1089), .A1(n960), .B0(N1276), .B1(n961), .Y(n959) );
  INVX1 U7660 ( .A(n962), .Y(n5795) );
  AOI22X1 U7661 ( .A0(N1088), .A1(n960), .B0(in_matrix_cnt[3]), .B1(n961), .Y(
        n962) );
  INVX1 U7662 ( .A(n963), .Y(n5794) );
  AOI22X1 U7663 ( .A0(N1087), .A1(n960), .B0(in_matrix_cnt[2]), .B1(n961), .Y(
        n963) );
  INVX1 U7664 ( .A(n964), .Y(n5793) );
  AOI22X1 U7665 ( .A0(N1086), .A1(n960), .B0(in_matrix_cnt[1]), .B1(n961), .Y(
        n964) );
  INVX1 U7666 ( .A(n965), .Y(n5792) );
  AOI22X1 U7667 ( .A0(N1085), .A1(n960), .B0(in_matrix_cnt[0]), .B1(n961), .Y(
        n965) );
  INVX1 U7668 ( .A(n958), .Y(n5798) );
  AOI21XL U7669 ( .A0(n925), .A1(in_weight_flag), .B0(N1276), .Y(n958) );
  AND2X2 U7670 ( .A(N1311), .B(n4474), .Y(N1321) );
  AND2X2 U7671 ( .A(N1339), .B(n5067), .Y(N1349) );
  AND3X2 U7672 ( .A(n1002), .B(n967), .C(in_valid), .Y(n994) );
  INVX1 U7673 ( .A(n993), .Y(n5824) );
  AOI22X1 U7674 ( .A0(n5832), .A1(in_cnt[7]), .B0(N1060), .B1(n994), .Y(n993)
         );
  NAND3X1 U7675 ( .A(in_cnt_64[1]), .B(in_cnt_64[0]), .C(in_cnt_64[2]), .Y(
        n1009) );
  NAND3X1 U7676 ( .A(in_cnt_64[4]), .B(in_cnt_64[3]), .C(in_cnt_64[5]), .Y(
        n1010) );
  NAND2X1 U7677 ( .A(n968), .B(in_valid), .Y(n4460) );
  AOI22X1 U7678 ( .A0(N1252), .A1(n5070), .B0(in_addr_cnt[9]), .B1(n5329), .Y(
        n968) );
  NAND2X1 U7679 ( .A(n971), .B(in_valid), .Y(n4461) );
  AOI22X1 U7680 ( .A0(N1251), .A1(n5070), .B0(n5329), .B1(in_addr_cnt[8]), .Y(
        n971) );
  NAND2X1 U7681 ( .A(n972), .B(in_valid), .Y(n4462) );
  AOI22X1 U7682 ( .A0(N1250), .A1(n5070), .B0(n5329), .B1(in_addr_cnt[7]), .Y(
        n972) );
  NAND2X1 U7683 ( .A(n973), .B(in_valid), .Y(n4463) );
  AOI22X1 U7684 ( .A0(N1249), .A1(n5070), .B0(n5329), .B1(in_addr_cnt[6]), .Y(
        n973) );
  NAND2X1 U7685 ( .A(n974), .B(in_valid), .Y(n4464) );
  AOI22X1 U7686 ( .A0(N1248), .A1(n5070), .B0(n5329), .B1(in_addr_cnt[5]), .Y(
        n974) );
  NAND2X1 U7687 ( .A(n975), .B(in_valid), .Y(n4465) );
  AOI22X1 U7688 ( .A0(N1247), .A1(n5070), .B0(n5329), .B1(in_addr_cnt[4]), .Y(
        n975) );
  NAND2X1 U7689 ( .A(n976), .B(in_valid), .Y(n4466) );
  AOI22X1 U7690 ( .A0(N1246), .A1(n5070), .B0(n5329), .B1(in_addr_cnt[3]), .Y(
        n976) );
  NAND2X1 U7691 ( .A(n977), .B(in_valid), .Y(n4467) );
  AOI22X1 U7692 ( .A0(N1245), .A1(n5070), .B0(n5329), .B1(in_addr_cnt[2]), .Y(
        n977) );
  NAND2X1 U7693 ( .A(n978), .B(in_valid), .Y(n4468) );
  AOI22X1 U7694 ( .A0(N1244), .A1(n5070), .B0(n5329), .B1(in_addr_cnt[1]), .Y(
        n978) );
  NAND2X1 U7695 ( .A(n979), .B(in_valid), .Y(n4469) );
  AOI22X1 U7696 ( .A0(N1243), .A1(n5070), .B0(n5329), .B1(in_addr_cnt[0]), .Y(
        n979) );
  NOR2BX1 U7697 ( .AN(in_valid), .B(n739), .Y(n970) );
  OAI2BB2X1 U7698 ( .B0(n1011), .B1(n5888), .A0N(matrix_size[1]), .A1N(n1011), 
        .Y(n4471) );
  OAI2BB2X1 U7699 ( .B0(n1011), .B1(n5886), .A0N(matrix_size[0]), .A1N(n1011), 
        .Y(n4470) );
  BUFX3 U7700 ( .A(n969), .Y(n5070) );
  AOI2BB1X1 U7701 ( .A0N(n980), .A1N(n981), .B0(n5329), .Y(n969) );
  NAND4X1 U7702 ( .A(in_addr_cnt[3]), .B(n989), .C(in_addr_cnt[2]), .D(n991), 
        .Y(n980) );
  NAND4X1 U7703 ( .A(n982), .B(n983), .C(n984), .D(n985), .Y(n981) );
  INVX1 U7704 ( .A(n995), .Y(n5825) );
  AOI22X1 U7705 ( .A0(n5832), .A1(in_cnt[6]), .B0(N1059), .B1(n994), .Y(n995)
         );
  INVX1 U7706 ( .A(n996), .Y(n5826) );
  AOI22X1 U7707 ( .A0(n5832), .A1(in_cnt[5]), .B0(N1058), .B1(n994), .Y(n996)
         );
  INVX1 U7708 ( .A(n997), .Y(n5827) );
  AOI22X1 U7709 ( .A0(n5832), .A1(in_cnt[4]), .B0(N1057), .B1(n994), .Y(n997)
         );
  INVX1 U7710 ( .A(n998), .Y(n5828) );
  AOI22X1 U7711 ( .A0(in_cnt[3]), .A1(n5832), .B0(N1056), .B1(n994), .Y(n998)
         );
  INVX1 U7712 ( .A(n999), .Y(n5829) );
  AOI22X1 U7713 ( .A0(in_cnt[2]), .A1(n5832), .B0(N1055), .B1(n994), .Y(n999)
         );
  INVX1 U7714 ( .A(n1000), .Y(n5830) );
  AOI22X1 U7715 ( .A0(in_cnt[1]), .A1(n5832), .B0(N1054), .B1(n994), .Y(n1000)
         );
  INVX1 U7716 ( .A(n1001), .Y(n5831) );
  AOI22X1 U7717 ( .A0(in_cnt[0]), .A1(n5832), .B0(N1053), .B1(n994), .Y(n1001)
         );
  AND2X2 U7718 ( .A(in_64[25]), .B(n5331), .Y(N1188) );
  AND2X2 U7719 ( .A(in_64[24]), .B(n5331), .Y(N1187) );
  AND2X2 U7720 ( .A(in_64[23]), .B(n5331), .Y(N1186) );
  AND2X2 U7721 ( .A(in_64[22]), .B(n5331), .Y(N1185) );
  AND2X2 U7722 ( .A(in_64[21]), .B(n5331), .Y(N1184) );
  AND2X2 U7723 ( .A(in_64[20]), .B(n5331), .Y(N1183) );
  AND2X2 U7724 ( .A(in_64[19]), .B(n5331), .Y(N1182) );
  AND2X2 U7725 ( .A(in_64[18]), .B(n5331), .Y(N1181) );
  AND2X2 U7726 ( .A(in_64[17]), .B(n5331), .Y(N1180) );
  AND2X2 U7727 ( .A(in_64[16]), .B(n5331), .Y(N1179) );
  AND2X2 U7728 ( .A(in_64[15]), .B(n5331), .Y(N1178) );
  AND2X2 U7729 ( .A(in_64[14]), .B(n5331), .Y(N1177) );
  AND2X2 U7730 ( .A(in_64[13]), .B(n5331), .Y(N1176) );
  AND2X2 U7731 ( .A(in_64[12]), .B(n5331), .Y(N1175) );
  AND2X2 U7732 ( .A(in_64[11]), .B(n5331), .Y(N1174) );
  AND2X2 U7733 ( .A(in_64[10]), .B(n5331), .Y(N1173) );
  AND2X2 U7734 ( .A(in_64[9]), .B(n5331), .Y(N1172) );
  AND2X2 U7735 ( .A(in_64[8]), .B(n5331), .Y(N1171) );
  AND2X2 U7736 ( .A(in_64[7]), .B(n5331), .Y(N1170) );
  AND2X2 U7737 ( .A(in_64[6]), .B(n5331), .Y(N1169) );
  AND2X2 U7738 ( .A(in_64[5]), .B(n5331), .Y(N1168) );
  AND2X2 U7739 ( .A(in_64[4]), .B(n5331), .Y(N1167) );
  AND2X2 U7740 ( .A(in_64[3]), .B(n5331), .Y(N1166) );
  AND2X2 U7741 ( .A(in_64[2]), .B(n5331), .Y(N1165) );
  AND2X2 U7742 ( .A(in_64[62]), .B(n5329), .Y(N1225) );
  AND2X2 U7743 ( .A(in_64[61]), .B(n5329), .Y(N1224) );
  AND2X2 U7744 ( .A(in_64[60]), .B(n5329), .Y(N1223) );
  AND2X2 U7745 ( .A(in_64[59]), .B(n5330), .Y(N1222) );
  AND2X2 U7746 ( .A(in_64[58]), .B(n5330), .Y(N1221) );
  AND2X2 U7747 ( .A(in_64[57]), .B(n5330), .Y(N1220) );
  AND2X2 U7748 ( .A(in_64[56]), .B(n5330), .Y(N1219) );
  AND2X2 U7749 ( .A(in_64[55]), .B(n5330), .Y(N1218) );
  AND2X2 U7750 ( .A(in_64[54]), .B(n5330), .Y(N1217) );
  AND2X2 U7751 ( .A(in_64[53]), .B(n5330), .Y(N1216) );
  AND2X2 U7752 ( .A(in_64[52]), .B(n5330), .Y(N1215) );
  AND2X2 U7753 ( .A(in_64[51]), .B(n5330), .Y(N1214) );
  AND2X2 U7754 ( .A(in_64[50]), .B(n5330), .Y(N1213) );
  AND2X2 U7755 ( .A(in_64[49]), .B(n5330), .Y(N1212) );
  AND2X2 U7756 ( .A(in_64[48]), .B(n5330), .Y(N1211) );
  AND2X2 U7757 ( .A(in_64[47]), .B(n5330), .Y(N1210) );
  AND2X2 U7758 ( .A(in_64[46]), .B(n5330), .Y(N1209) );
  AND2X2 U7759 ( .A(in_64[45]), .B(n5330), .Y(N1208) );
  AND2X2 U7760 ( .A(in_64[44]), .B(n5330), .Y(N1207) );
  AND2X2 U7761 ( .A(in_64[43]), .B(n5330), .Y(N1206) );
  AND2X2 U7762 ( .A(in_64[42]), .B(n5330), .Y(N1205) );
  AND2X2 U7763 ( .A(in_64[41]), .B(n5330), .Y(N1204) );
  AND2X2 U7764 ( .A(in_64[40]), .B(n5330), .Y(N1203) );
  AND2X2 U7765 ( .A(in_64[39]), .B(n5330), .Y(N1202) );
  AND2X2 U7766 ( .A(in_64[38]), .B(n5330), .Y(N1201) );
  AND2X2 U7767 ( .A(in_64[37]), .B(n5330), .Y(N1200) );
  AND2X2 U7768 ( .A(in_64[36]), .B(n5330), .Y(N1199) );
  AND2X2 U7769 ( .A(in_64[35]), .B(n5330), .Y(N1198) );
  AND2X2 U7770 ( .A(in_64[34]), .B(n5330), .Y(N1197) );
  AND2X2 U7771 ( .A(in_64[33]), .B(n5330), .Y(N1196) );
  AND2X2 U7772 ( .A(in_64[32]), .B(n5330), .Y(N1195) );
  AND2X2 U7773 ( .A(in_64[31]), .B(n5330), .Y(N1194) );
  AND2X2 U7774 ( .A(in_64[30]), .B(n5330), .Y(N1193) );
  AND2X2 U7775 ( .A(in_64[29]), .B(n5330), .Y(N1192) );
  AND2X2 U7776 ( .A(in_64[28]), .B(n5330), .Y(N1191) );
  AND2X2 U7777 ( .A(in_64[27]), .B(n5330), .Y(N1190) );
  AND2X2 U7778 ( .A(in_64[26]), .B(n5330), .Y(N1189) );
  AND2X2 U7779 ( .A(in_64[1]), .B(n5329), .Y(N1164) );
  AND2X2 U7780 ( .A(in_64[0]), .B(n5330), .Y(N1163) );
  NOR2BX1 U7781 ( .AN(w_mat[2]), .B(n5833), .Y(N1294) );
  NOR2BX1 U7782 ( .AN(w_mat[1]), .B(n5833), .Y(N1293) );
  NOR2BX1 U7783 ( .AN(w_mat[0]), .B(n5833), .Y(N1292) );
  NOR2BX1 U7784 ( .AN(w_mat_idx), .B(n5833), .Y(N1291) );
  NOR2BX1 U7785 ( .AN(i_mat[2]), .B(n5833), .Y(N1289) );
  NOR2BX1 U7786 ( .AN(i_mat[1]), .B(n5833), .Y(N1288) );
  NOR2BX1 U7787 ( .AN(i_mat[0]), .B(n5833), .Y(N1287) );
  NOR2BX1 U7788 ( .AN(i_mat_idx), .B(n5833), .Y(N1286) );
  AND2X2 U7789 ( .A(matrix), .B(in_valid), .Y(N1162) );
  AND2X2 U7790 ( .A(N1039), .B(in_valid), .Y(N1045) );
  AND2X2 U7791 ( .A(N1038), .B(in_valid), .Y(N1044) );
  AND2X2 U7792 ( .A(N1037), .B(in_valid), .Y(N1043) );
  AND2X2 U7793 ( .A(N1036), .B(in_valid), .Y(N1042) );
  AND2X2 U7794 ( .A(N1035), .B(in_valid), .Y(N1041) );
  AND2X2 U7795 ( .A(N1034), .B(in_valid), .Y(N1040) );
  CLKINVX3 U7796 ( .A(c_plus[34]), .Y(n5965) );
  NOR2X2 U7797 ( .A(cs[3]), .B(cs[0]), .Y(n1118) );
  OAI21X2 U7798 ( .A0(n5064), .A1(n5897), .B0(n1125), .Y(n1038) );
  OAI21XL U7799 ( .A0(store_cnt[3]), .A1(n5887), .B0(n1126), .Y(n1125) );
  OAI21XL U7800 ( .A0(n5885), .A1(n5896), .B0(n1127), .Y(n1126) );
  OAI21XL U7801 ( .A0(store_cnt[2]), .A1(n1128), .B0(n1129), .Y(n1127) );
  NAND3X1 U7802 ( .A(n851), .B(n787), .C(c_plus[14]), .Y(n815) );
  NAND2X1 U7803 ( .A(m_size[1]), .B(n5887), .Y(n1045) );
  INVX4 U7804 ( .A(c_plus[35]), .Y(n5966) );
  CLKINVX3 U7805 ( .A(cs[1]), .Y(n5890) );
  INVX1 U7806 ( .A(m_size[1]), .Y(n5888) );
  NAND4X1 U7807 ( .A(n812), .B(n793), .C(n815), .D(n850), .Y(n833) );
  AOI22X1 U7808 ( .A0(c_plus[6]), .A1(n832), .B0(c_plus[38]), .B1(n5970), .Y(
        n850) );
  BUFX3 U7809 ( .A(n761), .Y(n5080) );
  NOR4BX1 U7810 ( .AN(n825), .B(n820), .C(n826), .D(n827), .Y(n761) );
  NAND4X1 U7811 ( .A(c_plus[1]), .B(n819), .C(n5966), .D(n5933), .Y(n825) );
  NAND4X1 U7812 ( .A(n785), .B(n805), .C(n799), .D(n778), .Y(n827) );
  BUFX3 U7813 ( .A(n690), .Y(n5085) );
  BUFX3 U7814 ( .A(n760), .Y(n5081) );
  AND4X2 U7815 ( .A(n809), .B(n790), .C(n817), .D(n818), .Y(n760) );
  AOI21X1 U7816 ( .A0(c_plus[35]), .A1(n5970), .B0(n796), .Y(n817) );
  AOI211X1 U7817 ( .A0(c_plus[3]), .A1(n819), .B0(n820), .C0(n821), .Y(n818)
         );
  OAI2BB2X1 U7818 ( .B0(n5081), .B1(n5637), .A0N(length_reg[86]), .A1N(n5857), 
        .Y(n1725) );
  OAI2BB2X1 U7819 ( .B0(n5080), .B1(n5636), .A0N(length_reg[85]), .A1N(n5857), 
        .Y(n1726) );
  OAI2BB2X1 U7820 ( .B0(n5081), .B1(n5594), .A0N(length_reg[2]), .A1N(n5191), 
        .Y(n1809) );
  OAI2BB2X1 U7821 ( .B0(n5081), .B1(n5597), .A0N(length_reg[8]), .A1N(n5195), 
        .Y(n1803) );
  OAI2BB2X1 U7822 ( .B0(n5081), .B1(n5600), .A0N(length_reg[14]), .A1N(n5199), 
        .Y(n1797) );
  OAI2BB2X1 U7823 ( .B0(n5081), .B1(n5603), .A0N(length_reg[20]), .A1N(n5203), 
        .Y(n1791) );
  OAI2BB2X1 U7824 ( .B0(n5081), .B1(n5606), .A0N(length_reg[26]), .A1N(n5207), 
        .Y(n1785) );
  OAI2BB2X1 U7825 ( .B0(n5081), .B1(n5609), .A0N(length_reg[32]), .A1N(n5211), 
        .Y(n1779) );
  OAI2BB2X1 U7826 ( .B0(n5081), .B1(n5612), .A0N(length_reg[38]), .A1N(n5215), 
        .Y(n1773) );
  OAI2BB2X1 U7827 ( .B0(n5081), .B1(n5615), .A0N(length_reg[44]), .A1N(n5219), 
        .Y(n1767) );
  OAI2BB2X1 U7828 ( .B0(n5081), .B1(n5618), .A0N(length_reg[50]), .A1N(n5223), 
        .Y(n1761) );
  OAI2BB2X1 U7829 ( .B0(n5081), .B1(n5621), .A0N(length_reg[56]), .A1N(n5227), 
        .Y(n1755) );
  OAI2BB2X1 U7830 ( .B0(n5081), .B1(n5624), .A0N(length_reg[62]), .A1N(n5231), 
        .Y(n1749) );
  OAI2BB2X1 U7831 ( .B0(n5081), .B1(n5627), .A0N(length_reg[68]), .A1N(n5233), 
        .Y(n1743) );
  OAI2BB2X1 U7832 ( .B0(n5081), .B1(n5630), .A0N(length_reg[74]), .A1N(n5239), 
        .Y(n1737) );
  OAI2BB2X1 U7833 ( .B0(n5081), .B1(n5633), .A0N(length_reg[80]), .A1N(n5243), 
        .Y(n1731) );
  OAI2BB2X1 U7834 ( .B0(n5080), .B1(n5594), .A0N(length_reg[1]), .A1N(n5843), 
        .Y(n1810) );
  OAI2BB2X1 U7835 ( .B0(n5080), .B1(n5597), .A0N(length_reg[7]), .A1N(n5844), 
        .Y(n1804) );
  OAI2BB2X1 U7836 ( .B0(n5080), .B1(n5600), .A0N(length_reg[13]), .A1N(n5845), 
        .Y(n1798) );
  OAI2BB2X1 U7837 ( .B0(n5080), .B1(n5603), .A0N(length_reg[19]), .A1N(n5846), 
        .Y(n1792) );
  OAI2BB2X1 U7838 ( .B0(n5080), .B1(n5606), .A0N(length_reg[25]), .A1N(n5847), 
        .Y(n1786) );
  OAI2BB2X1 U7839 ( .B0(n5080), .B1(n5609), .A0N(length_reg[31]), .A1N(n5848), 
        .Y(n1780) );
  OAI2BB2X1 U7840 ( .B0(n5080), .B1(n5612), .A0N(length_reg[37]), .A1N(n5849), 
        .Y(n1774) );
  OAI2BB2X1 U7841 ( .B0(n5080), .B1(n5615), .A0N(length_reg[43]), .A1N(n5850), 
        .Y(n1768) );
  OAI2BB2X1 U7842 ( .B0(n5080), .B1(n5618), .A0N(length_reg[49]), .A1N(n5851), 
        .Y(n1762) );
  OAI2BB2X1 U7843 ( .B0(n5080), .B1(n5621), .A0N(length_reg[55]), .A1N(n5852), 
        .Y(n1756) );
  OAI2BB2X1 U7844 ( .B0(n5080), .B1(n5624), .A0N(length_reg[61]), .A1N(n5853), 
        .Y(n1750) );
  OAI2BB2X1 U7845 ( .B0(n5080), .B1(n5627), .A0N(length_reg[67]), .A1N(n5854), 
        .Y(n1744) );
  OAI2BB2X1 U7846 ( .B0(n5080), .B1(n5630), .A0N(length_reg[73]), .A1N(n5855), 
        .Y(n1738) );
  OAI2BB2X1 U7847 ( .B0(n5080), .B1(n5633), .A0N(length_reg[79]), .A1N(n5243), 
        .Y(n1732) );
  NAND4X1 U7848 ( .A(n811), .B(n792), .C(n816), .D(n831), .Y(n820) );
  BUFX3 U7849 ( .A(mem_num_4_), .Y(n5064) );
  NOR2X1 U7850 ( .A(n5888), .B(m_size[0]), .Y(mem_num_4_) );
  NAND4X1 U7851 ( .A(n794), .B(n781), .C(n810), .D(n855), .Y(n821) );
  AOI31X1 U7852 ( .A0(n832), .A1(n5935), .A2(c_plus[4]), .B0(n795), .Y(n855)
         );
  NOR2X2 U7853 ( .A(out_cnt[0]), .B(out_cnt[1]), .Y(n1059) );
  NAND4X1 U7854 ( .A(n1040), .B(n4890), .C(n1041), .D(n1042), .Y(n1039) );
  XNOR2X1 U7855 ( .A(N944), .B(n5885), .Y(n1041) );
  XNOR2X1 U7856 ( .A(N943), .B(n1045), .Y(n1040) );
  CLKINVX3 U7857 ( .A(c_plus[19]), .Y(n5950) );
  CLKINVX3 U7858 ( .A(c_plus[18]), .Y(n5949) );
  CLKINVX3 U7859 ( .A(c_plus[28]), .Y(n5960) );
  CLKINVX3 U7860 ( .A(c_plus[23]), .Y(n5954) );
  CLKINVX3 U7861 ( .A(c_plus[27]), .Y(n5959) );
  AND4X2 U7862 ( .A(n5250), .B(n4492), .C(n4493), .D(n4494), .Y(n1132) );
  XOR2X1 U7863 ( .A(n1128), .B(calin_cnt[0]), .Y(n4492) );
  XOR2X1 U7864 ( .A(calin_cnt[3]), .B(n5887), .Y(n4493) );
  XOR2X1 U7865 ( .A(calin_cnt[2]), .B(n5887), .Y(n4494) );
  NAND3X1 U7866 ( .A(n822), .B(n5942), .C(c_plus[10]), .Y(n800) );
  INVX1 U7867 ( .A(n1030), .Y(n5834) );
  AOI22X1 U7868 ( .A0(N14363), .A1(n1031), .B0(N14369), .B1(n1032), .Y(n1030)
         );
  AOI31X1 U7869 ( .A0(c_plus[2]), .A1(n832), .A2(n853), .B0(n5941), .Y(n852)
         );
  NOR3X1 U7870 ( .A(c_plus[3]), .B(c_plus[5]), .C(c_plus[4]), .Y(n853) );
  INVX1 U7871 ( .A(n800), .Y(n5941) );
  AOI22X1 U7872 ( .A0(value_out[4]), .A1(n1059), .B0(value_out[7]), .B1(n1060), 
        .Y(n1079) );
  AOI22X1 U7873 ( .A0(value_out[12]), .A1(n1059), .B0(value_out[15]), .B1(
        n1060), .Y(n1074) );
  AOI22X1 U7874 ( .A0(value_out[20]), .A1(n1059), .B0(value_out[23]), .B1(
        n1060), .Y(n1058) );
  AOI22X1 U7875 ( .A0(value_out[36]), .A1(n1059), .B0(value_out[39]), .B1(
        n1060), .Y(n1084) );
  AOI22X1 U7876 ( .A0(value_out[6]), .A1(n1061), .B0(value_out[5]), .B1(n1062), 
        .Y(n1078) );
  AOI22X1 U7877 ( .A0(value_out[14]), .A1(n1061), .B0(value_out[13]), .B1(
        n1062), .Y(n1073) );
  AOI22X1 U7878 ( .A0(value_out[22]), .A1(n1061), .B0(value_out[21]), .B1(
        n1062), .Y(n1057) );
  AOI22X1 U7879 ( .A0(value_out[38]), .A1(n1061), .B0(value_out[37]), .B1(
        n1062), .Y(n1083) );
  AOI22X1 U7880 ( .A0(n1051), .A1(n5976), .B0(out_cnt[4]), .B1(n1052), .Y(
        n1050) );
  OAI22X1 U7881 ( .A0(n1053), .A1(n5975), .B0(out_cnt[3]), .B1(n1054), .Y(
        n1052) );
  OAI32X1 U7882 ( .A0(n1069), .A1(out_cnt[5]), .A2(out_cnt[3]), .B0(n1070), 
        .B1(n5975), .Y(n1051) );
  AOI211X1 U7883 ( .A0(value_out[24]), .A1(n1044), .B0(n1064), .C0(n1065), .Y(
        n1053) );
  AOI22X1 U7884 ( .A0(calin_cnt[3]), .A1(n5061), .B0(n5064), .B1(calin_cnt[4]), 
        .Y(n955) );
  NAND3X1 U7885 ( .A(n787), .B(n5948), .C(c_plus[16]), .Y(n784) );
  NAND3X1 U7886 ( .A(n836), .B(n5952), .C(c_plus[20]), .Y(n794) );
  NAND3X1 U7887 ( .A(n823), .B(n5950), .C(c_plus[18]), .Y(n791) );
  NAND2X1 U7888 ( .A(c_plus[24]), .B(n813), .Y(n814) );
  NAND3X1 U7889 ( .A(cs[1]), .B(n1118), .C(cs[2]), .Y(n1120) );
  NOR2BX1 U7890 ( .AN(calin_cnt[0]), .B(n5887), .Y(n956) );
  AND4X2 U7891 ( .A(n5949), .B(n5950), .C(n851), .D(n857), .Y(n834) );
  NOR3X1 U7892 ( .A(c_plus[20]), .B(c_plus[22]), .C(c_plus[21]), .Y(n857) );
  NAND2X1 U7893 ( .A(c_plus[22]), .B(n835), .Y(n793) );
  INVX1 U7894 ( .A(m_size[0]), .Y(n5886) );
  NOR2X1 U7895 ( .A(out_cnt[2]), .B(n1068), .Y(n1064) );
  AOI211X1 U7896 ( .A0(value_out[32]), .A1(n1044), .B0(n1081), .C0(n1082), .Y(
        n1049) );
  AOI21X1 U7897 ( .A0(n1083), .A1(n1084), .B0(n5974), .Y(n1082) );
  NOR2X1 U7898 ( .A(out_cnt[2]), .B(n1085), .Y(n1081) );
  BUFX3 U7899 ( .A(n1014), .Y(n5066) );
  NAND3X1 U7900 ( .A(n1118), .B(n5889), .C(cs[1]), .Y(n1014) );
  NOR2X1 U7901 ( .A(n1046), .B(n746), .Y(N14331) );
  AOI22X1 U7902 ( .A0(n1047), .A1(n5973), .B0(n1012), .B1(n1048), .Y(n1046) );
  OAI22X1 U7903 ( .A0(n1086), .A1(n728), .B0(out_cnt_6[0]), .B1(n1087), .Y(
        n1047) );
  OAI21XL U7904 ( .A0(n1049), .A1(n5977), .B0(n1050), .Y(n1048) );
  NAND2X1 U7905 ( .A(c_plus[17]), .B(n787), .Y(n785) );
  NAND2X1 U7906 ( .A(c_plus[21]), .B(n836), .Y(n792) );
  BUFX3 U7907 ( .A(n758), .Y(n5083) );
  AND4X2 U7908 ( .A(n783), .B(n784), .C(n785), .D(n786), .Y(n758) );
  AND3X2 U7909 ( .A(n789), .B(n790), .C(n791), .Y(n783) );
  AOI21X1 U7910 ( .A0(c_plus[15]), .A1(n787), .B0(n788), .Y(n786) );
  OAI2BB2X1 U7911 ( .B0(n5079), .B1(n5636), .A0N(length_reg[84]), .A1N(n5857), 
        .Y(n1727) );
  OAI2BB2X1 U7912 ( .B0(n5083), .B1(n5637), .A0N(length_reg[88]), .A1N(n5857), 
        .Y(n1723) );
  OAI2BB2X1 U7913 ( .B0(n5082), .B1(n5637), .A0N(length_reg[87]), .A1N(n5857), 
        .Y(n1724) );
  AND2X2 U7914 ( .A(n822), .B(c_plus[11]), .Y(n796) );
  OAI2BB2X1 U7915 ( .B0(n5079), .B1(n5594), .A0N(length_reg[0]), .A1N(n5843), 
        .Y(n1811) );
  OAI2BB2X1 U7916 ( .B0(n5079), .B1(n5597), .A0N(length_reg[6]), .A1N(n5844), 
        .Y(n1805) );
  OAI2BB2X1 U7917 ( .B0(n5079), .B1(n5600), .A0N(length_reg[12]), .A1N(n5845), 
        .Y(n1799) );
  OAI2BB2X1 U7918 ( .B0(n5079), .B1(n5603), .A0N(length_reg[18]), .A1N(n5846), 
        .Y(n1793) );
  OAI2BB2X1 U7919 ( .B0(n5079), .B1(n5606), .A0N(length_reg[24]), .A1N(n5847), 
        .Y(n1787) );
  OAI2BB2X1 U7920 ( .B0(n5079), .B1(n5609), .A0N(length_reg[30]), .A1N(n5848), 
        .Y(n1781) );
  OAI2BB2X1 U7921 ( .B0(n5079), .B1(n5612), .A0N(length_reg[36]), .A1N(n5849), 
        .Y(n1775) );
  OAI2BB2X1 U7922 ( .B0(n5079), .B1(n5615), .A0N(length_reg[42]), .A1N(n5850), 
        .Y(n1769) );
  OAI2BB2X1 U7923 ( .B0(n5079), .B1(n5618), .A0N(length_reg[48]), .A1N(n5851), 
        .Y(n1763) );
  OAI2BB2X1 U7924 ( .B0(n5079), .B1(n5621), .A0N(length_reg[54]), .A1N(n5852), 
        .Y(n1757) );
  OAI2BB2X1 U7925 ( .B0(n5079), .B1(n5624), .A0N(length_reg[60]), .A1N(n5853), 
        .Y(n1751) );
  OAI2BB2X1 U7926 ( .B0(n5079), .B1(n5627), .A0N(length_reg[66]), .A1N(n5854), 
        .Y(n1745) );
  OAI2BB2X1 U7927 ( .B0(n5079), .B1(n5630), .A0N(length_reg[72]), .A1N(n5855), 
        .Y(n1739) );
  OAI2BB2X1 U7928 ( .B0(n5079), .B1(n5633), .A0N(length_reg[78]), .A1N(n5243), 
        .Y(n1733) );
  OAI2BB2X1 U7929 ( .B0(n5083), .B1(n5594), .A0N(length_reg[4]), .A1N(n5843), 
        .Y(n1807) );
  OAI2BB2X1 U7930 ( .B0(n5083), .B1(n5597), .A0N(length_reg[10]), .A1N(n5844), 
        .Y(n1801) );
  OAI2BB2X1 U7931 ( .B0(n5083), .B1(n5600), .A0N(length_reg[16]), .A1N(n5845), 
        .Y(n1795) );
  OAI2BB2X1 U7932 ( .B0(n5083), .B1(n5603), .A0N(length_reg[22]), .A1N(n5846), 
        .Y(n1789) );
  OAI2BB2X1 U7933 ( .B0(n5083), .B1(n5606), .A0N(length_reg[28]), .A1N(n5847), 
        .Y(n1783) );
  OAI2BB2X1 U7934 ( .B0(n5083), .B1(n5609), .A0N(length_reg[34]), .A1N(n5848), 
        .Y(n1777) );
  OAI2BB2X1 U7935 ( .B0(n5083), .B1(n5612), .A0N(length_reg[40]), .A1N(n5849), 
        .Y(n1771) );
  OAI2BB2X1 U7936 ( .B0(n5083), .B1(n5615), .A0N(length_reg[46]), .A1N(n5850), 
        .Y(n1765) );
  OAI2BB2X1 U7937 ( .B0(n5083), .B1(n5618), .A0N(length_reg[52]), .A1N(n5851), 
        .Y(n1759) );
  OAI2BB2X1 U7938 ( .B0(n5083), .B1(n5621), .A0N(length_reg[58]), .A1N(n5852), 
        .Y(n1753) );
  OAI2BB2X1 U7939 ( .B0(n5083), .B1(n5624), .A0N(length_reg[64]), .A1N(n5853), 
        .Y(n1747) );
  OAI2BB2X1 U7940 ( .B0(n5083), .B1(n5627), .A0N(length_reg[70]), .A1N(n5854), 
        .Y(n1741) );
  OAI2BB2X1 U7941 ( .B0(n5083), .B1(n5630), .A0N(length_reg[76]), .A1N(n5855), 
        .Y(n1735) );
  OAI2BB2X1 U7942 ( .B0(n5083), .B1(n5633), .A0N(length_reg[82]), .A1N(n5243), 
        .Y(n1729) );
  OAI2BB2X1 U7943 ( .B0(n5082), .B1(n5594), .A0N(length_reg[3]), .A1N(n5843), 
        .Y(n1808) );
  OAI2BB2X1 U7944 ( .B0(n5082), .B1(n5597), .A0N(length_reg[9]), .A1N(n5844), 
        .Y(n1802) );
  OAI2BB2X1 U7945 ( .B0(n5082), .B1(n5600), .A0N(length_reg[15]), .A1N(n5845), 
        .Y(n1796) );
  OAI2BB2X1 U7946 ( .B0(n5082), .B1(n5603), .A0N(length_reg[21]), .A1N(n5846), 
        .Y(n1790) );
  OAI2BB2X1 U7947 ( .B0(n5082), .B1(n5606), .A0N(length_reg[27]), .A1N(n5847), 
        .Y(n1784) );
  OAI2BB2X1 U7948 ( .B0(n5082), .B1(n5609), .A0N(length_reg[33]), .A1N(n5848), 
        .Y(n1778) );
  OAI2BB2X1 U7949 ( .B0(n5082), .B1(n5612), .A0N(length_reg[39]), .A1N(n5849), 
        .Y(n1772) );
  OAI2BB2X1 U7950 ( .B0(n5082), .B1(n5615), .A0N(length_reg[45]), .A1N(n5850), 
        .Y(n1766) );
  OAI2BB2X1 U7951 ( .B0(n5082), .B1(n5618), .A0N(length_reg[51]), .A1N(n5851), 
        .Y(n1760) );
  OAI2BB2X1 U7952 ( .B0(n5082), .B1(n5621), .A0N(length_reg[57]), .A1N(n5852), 
        .Y(n1754) );
  OAI2BB2X1 U7953 ( .B0(n5082), .B1(n5624), .A0N(length_reg[63]), .A1N(n5853), 
        .Y(n1748) );
  OAI2BB2X1 U7954 ( .B0(n5082), .B1(n5627), .A0N(length_reg[69]), .A1N(n5854), 
        .Y(n1742) );
  OAI2BB2X1 U7955 ( .B0(n5082), .B1(n5630), .A0N(length_reg[75]), .A1N(n5855), 
        .Y(n1736) );
  OAI2BB2X1 U7956 ( .B0(n5082), .B1(n5633), .A0N(length_reg[81]), .A1N(n5243), 
        .Y(n1730) );
  NAND2X1 U7957 ( .A(c_plus[19]), .B(n823), .Y(n790) );
  AOI211X1 U7958 ( .A0(value_out[16]), .A1(n1044), .B0(n1055), .C0(n1056), .Y(
        n1054) );
  AOI21X1 U7959 ( .A0(n1057), .A1(n1058), .B0(n5974), .Y(n1056) );
  NOR2X1 U7960 ( .A(out_cnt[2]), .B(n1063), .Y(n1055) );
  INVX1 U7961 ( .A(N944), .Y(n4889) );
  XNOR2X1 U7962 ( .A(calin_cnt[1]), .B(n5885), .Y(n1130) );
  INVX1 U7963 ( .A(N942), .Y(n4890) );
  AOI31X1 U7964 ( .A0(c_plus[7]), .A1(n803), .A2(n804), .B0(n788), .Y(n802) );
  NOR3X1 U7965 ( .A(c_plus[35]), .B(c_plus[38]), .C(c_plus[37]), .Y(n804) );
  BUFX3 U7966 ( .A(mem_num_2), .Y(n5061) );
  NOR2X1 U7967 ( .A(n5886), .B(m_size[1]), .Y(mem_num_2) );
  AND2X2 U7968 ( .A(n856), .B(c_plus[12]), .Y(n795) );
  INVX1 U7969 ( .A(n1033), .Y(n5835) );
  AOI22X1 U7970 ( .A0(N14362), .A1(n1031), .B0(N14368), .B1(n1032), .Y(n1033)
         );
  INVX1 U7971 ( .A(n1034), .Y(n5836) );
  AOI22X1 U7972 ( .A0(N14361), .A1(n1031), .B0(N14367), .B1(n1032), .Y(n1034)
         );
  XNOR2X1 U7973 ( .A(N945), .B(n5887), .Y(n1043) );
  NAND4X1 U7974 ( .A(n805), .B(n806), .C(n807), .D(n808), .Y(n788) );
  AND4X2 U7975 ( .A(n809), .B(n810), .C(n811), .D(n812), .Y(n808) );
  AOI21X1 U7976 ( .A0(c_plus[23]), .A1(n813), .B0(n5956), .Y(n807) );
  INVX1 U7977 ( .A(n814), .Y(n5956) );
  AOI211X1 U7978 ( .A0(value_out[0]), .A1(n1044), .B0(n1076), .C0(n1077), .Y(
        n1069) );
  AOI21X1 U7979 ( .A0(n1078), .A1(n1079), .B0(n5974), .Y(n1077) );
  NOR2X1 U7980 ( .A(out_cnt[2]), .B(n1080), .Y(n1076) );
  AOI211X1 U7981 ( .A0(value_out[8]), .A1(n1044), .B0(n1071), .C0(n1072), .Y(
        n1070) );
  AOI21X1 U7982 ( .A0(n1073), .A1(n1074), .B0(n5974), .Y(n1072) );
  NOR2X1 U7983 ( .A(out_cnt[2]), .B(n1075), .Y(n1071) );
  CLKINVX3 U7984 ( .A(c_plus[22]), .Y(n5953) );
  CLKINVX3 U7985 ( .A(c_plus[7]), .Y(n5937) );
  CLKINVX3 U7986 ( .A(c_plus[13]), .Y(n5944) );
  CLKINVX3 U7987 ( .A(c_plus[20]), .Y(n5951) );
  AND4X2 U7988 ( .A(n966), .B(in_cnt_64[4]), .C(in_cnt_64[3]), .D(in_cnt_64[5]), .Y(n960) );
  AND4X2 U7989 ( .A(n5884), .B(in_cnt_64[0]), .C(in_cnt_64[1]), .D(
        in_cnt_64[2]), .Y(n966) );
  INVX1 U7990 ( .A(n967), .Y(n5884) );
  AND2X2 U7991 ( .A(out_cnt[1]), .B(n5971), .Y(n1061) );
  AND2X2 U7992 ( .A(out_cnt[1]), .B(out_cnt[0]), .Y(n1060) );
  INVX1 U7993 ( .A(n1036), .Y(n5838) );
  AOI22X1 U7994 ( .A0(N14359), .A1(n1031), .B0(N14365), .B1(n1032), .Y(n1036)
         );
  INVX1 U7995 ( .A(n1037), .Y(n5839) );
  AOI22XL U7996 ( .A0(N14358), .A1(n1031), .B0(n5971), .B1(n1032), .Y(n1037)
         );
  OR2X2 U7997 ( .A(r1350_GE_LT_GT_LE), .B(n5050), .Y(n1649) );
  INVX1 U7998 ( .A(n5649), .Y(n5654) );
  INVXL U7999 ( .A(mem_num_0), .Y(n5662) );
  INVX4 U8000 ( .A(c_plus[39]), .Y(n5970) );
  NOR4X1 U8001 ( .A(in_cnt[7]), .B(in_cnt[6]), .C(in_cnt[5]), .D(in_cnt[4]), 
        .Y(n1006) );
  XNOR2X1 U8002 ( .A(in_cnt[0]), .B(n5885), .Y(n1003) );
  XNOR2X1 U8003 ( .A(in_cnt[1]), .B(n5885), .Y(n1004) );
  OAI22X1 U8004 ( .A0(n465), .A1(n5309), .B0(n497), .B1(n5263), .Y(n1317) );
  OAI22X1 U8005 ( .A0(n609), .A1(n5310), .B0(n657), .B1(n5261), .Y(n1582) );
  OAI22X1 U8006 ( .A0(n464), .A1(n5310), .B0(n496), .B1(n5263), .Y(n1313) );
  OAI22X1 U8007 ( .A0(n608), .A1(n5310), .B0(n656), .B1(n5261), .Y(n1578) );
  OAI22X1 U8008 ( .A0(n463), .A1(n5309), .B0(n495), .B1(n5263), .Y(n1309) );
  OAI22X1 U8009 ( .A0(n607), .A1(n5309), .B0(n655), .B1(n5261), .Y(n1574) );
  OAI22X1 U8010 ( .A0(n462), .A1(n5310), .B0(n494), .B1(n5263), .Y(n1305) );
  OAI22X1 U8011 ( .A0(n606), .A1(n5310), .B0(n654), .B1(n5261), .Y(n1570) );
  OAI22X1 U8012 ( .A0(n461), .A1(n5310), .B0(n493), .B1(n5263), .Y(n1301) );
  OAI22X1 U8013 ( .A0(n605), .A1(n5309), .B0(n653), .B1(n5261), .Y(n1566) );
  OAI22X1 U8014 ( .A0(n460), .A1(n5310), .B0(n492), .B1(n5263), .Y(n1297) );
  OAI22X1 U8015 ( .A0(n604), .A1(n5310), .B0(n652), .B1(n5261), .Y(n1562) );
  OAI22X1 U8016 ( .A0(n459), .A1(n5310), .B0(n491), .B1(n5263), .Y(n1293) );
  OAI22X1 U8017 ( .A0(n603), .A1(n5309), .B0(n651), .B1(n5261), .Y(n1558) );
  OAI22X1 U8018 ( .A0(n602), .A1(n5309), .B0(n650), .B1(n5261), .Y(n1554) );
  OAI22X1 U8019 ( .A0(n601), .A1(n5309), .B0(n649), .B1(n5261), .Y(n1550) );
  OAI22X1 U8020 ( .A0(n600), .A1(n5309), .B0(n648), .B1(n5261), .Y(n1546) );
  OAI22X1 U8021 ( .A0(n599), .A1(n5308), .B0(n647), .B1(n5261), .Y(n1542) );
  OAI22X1 U8022 ( .A0(n598), .A1(n5310), .B0(n646), .B1(n5261), .Y(n1538) );
  OAI22X1 U8023 ( .A0(n597), .A1(n5308), .B0(n645), .B1(n5261), .Y(n1534) );
  OAI22X1 U8024 ( .A0(n596), .A1(n5309), .B0(n644), .B1(n5262), .Y(n1530) );
  OAI22X1 U8025 ( .A0(n595), .A1(n5308), .B0(n643), .B1(n5262), .Y(n1526) );
  OAI22X1 U8026 ( .A0(n594), .A1(n5309), .B0(n642), .B1(n5262), .Y(n1521) );
  OAI22X1 U8027 ( .A0(n529), .A1(n5307), .B0(n561), .B1(n5262), .Y(n1449) );
  OAI22X1 U8028 ( .A0(n528), .A1(n5308), .B0(n560), .B1(n5262), .Y(n1445) );
  OAI22X1 U8029 ( .A0(n527), .A1(n5308), .B0(n559), .B1(n5262), .Y(n1441) );
  OAI22X1 U8030 ( .A0(n526), .A1(n5309), .B0(n558), .B1(n5262), .Y(n1437) );
  OAI22X1 U8031 ( .A0(n525), .A1(n5308), .B0(n557), .B1(n5262), .Y(n1433) );
  OAI22X1 U8032 ( .A0(n524), .A1(n5308), .B0(n556), .B1(n5262), .Y(n1429) );
  OAI22X1 U8033 ( .A0(n523), .A1(n5308), .B0(n555), .B1(n5262), .Y(n1425) );
  OAI22X1 U8034 ( .A0(n522), .A1(n5310), .B0(n554), .B1(n5262), .Y(n1421) );
  OAI22X1 U8035 ( .A0(n521), .A1(n5308), .B0(n553), .B1(n5262), .Y(n1417) );
  OAI22X1 U8036 ( .A0(n520), .A1(n5309), .B0(n552), .B1(n5262), .Y(n1413) );
  OAI22X1 U8037 ( .A0(n519), .A1(n5308), .B0(n551), .B1(n5263), .Y(n1409) );
  OAI22X1 U8038 ( .A0(n518), .A1(n5308), .B0(n550), .B1(n5263), .Y(n1405) );
  OAI22X1 U8039 ( .A0(n517), .A1(n5308), .B0(n549), .B1(n5263), .Y(n1401) );
  OAI22X1 U8040 ( .A0(n516), .A1(n5309), .B0(n548), .B1(n5263), .Y(n1397) );
  OAI22X1 U8041 ( .A0(n515), .A1(n5308), .B0(n547), .B1(n5263), .Y(n1393) );
  OAI22X1 U8042 ( .A0(n514), .A1(n5310), .B0(n546), .B1(n5263), .Y(n1388) );
  OAI22X1 U8043 ( .A0(n593), .A1(n5284), .B0(n641), .B1(n5304), .Y(n1650) );
  OAI22X1 U8044 ( .A0(n375), .A1(n5286), .B0(n423), .B1(n5304), .Y(n1209) );
  OAI22X1 U8045 ( .A0(n374), .A1(n5285), .B0(n422), .B1(n5304), .Y(n1205) );
  OAI22X1 U8046 ( .A0(n582), .A1(n5284), .B0(n630), .B1(n5307), .Y(n1604) );
  OAI22X1 U8047 ( .A0(n373), .A1(n5285), .B0(n421), .B1(n5304), .Y(n1201) );
  OAI22X1 U8048 ( .A0(n372), .A1(n5285), .B0(n420), .B1(n5304), .Y(n1197) );
  OAI22X1 U8049 ( .A0(n371), .A1(n5284), .B0(n419), .B1(n5304), .Y(n1193) );
  OAI22X1 U8050 ( .A0(n590), .A1(n5284), .B0(n638), .B1(n5307), .Y(n1636) );
  OAI22X1 U8051 ( .A0(n589), .A1(n5284), .B0(n637), .B1(n5307), .Y(n1632) );
  OAI22X1 U8052 ( .A0(n588), .A1(n5284), .B0(n636), .B1(n5307), .Y(n1628) );
  OAI22X1 U8053 ( .A0(n382), .A1(n5287), .B0(n430), .B1(n5304), .Y(n1237) );
  OAI22X1 U8054 ( .A0(n381), .A1(n5287), .B0(n429), .B1(n5304), .Y(n1233) );
  OAI22X1 U8055 ( .A0(n380), .A1(n5284), .B0(n428), .B1(n5304), .Y(n1229) );
  OAI22X1 U8056 ( .A0(n379), .A1(n5287), .B0(n427), .B1(n5304), .Y(n1225) );
  OAI22X1 U8057 ( .A0(n378), .A1(n5284), .B0(n426), .B1(n5304), .Y(n1221) );
  OAI22X1 U8058 ( .A0(n377), .A1(n5287), .B0(n425), .B1(n5304), .Y(n1217) );
  OAI22X1 U8059 ( .A0(n376), .A1(n5286), .B0(n424), .B1(n5304), .Y(n1213) );
  OAI22X1 U8060 ( .A0(n385), .A1(n5287), .B0(n433), .B1(n5305), .Y(n1249) );
  OAI22X1 U8061 ( .A0(n513), .A1(n5285), .B0(n545), .B1(n5307), .Y(n1515) );
  OAI22X1 U8062 ( .A0(n503), .A1(n5286), .B0(n535), .B1(n5306), .Y(n1475) );
  OAI22X1 U8063 ( .A0(n583), .A1(n5284), .B0(n631), .B1(n5307), .Y(n1608) );
  OAI22X1 U8064 ( .A0(n502), .A1(n5286), .B0(n534), .B1(n5307), .Y(n1471) );
  OAI22X1 U8065 ( .A0(n501), .A1(n5286), .B0(n533), .B1(n5306), .Y(n1467) );
  OAI22X1 U8066 ( .A0(n581), .A1(n5284), .B0(n629), .B1(n5307), .Y(n1600) );
  OAI22X1 U8067 ( .A0(n500), .A1(n5286), .B0(n532), .B1(n5307), .Y(n1463) );
  OAI22X1 U8068 ( .A0(n580), .A1(n5285), .B0(n628), .B1(n5306), .Y(n1596) );
  OAI22X1 U8069 ( .A0(n499), .A1(n5286), .B0(n531), .B1(n5306), .Y(n1459) );
  OAI22X1 U8070 ( .A0(n579), .A1(n5285), .B0(n627), .B1(n5307), .Y(n1592) );
  OAI22X1 U8071 ( .A0(n370), .A1(n5297), .B0(n418), .B1(n5305), .Y(n1184) );
  OAI22X1 U8072 ( .A0(n498), .A1(n5286), .B0(n530), .B1(n5307), .Y(n1454) );
  OAI22X1 U8073 ( .A0(n578), .A1(n5285), .B0(n626), .B1(n5306), .Y(n1587) );
  OAI22X1 U8074 ( .A0(n384), .A1(n5287), .B0(n432), .B1(n5306), .Y(n1245) );
  OAI22X1 U8075 ( .A0(n512), .A1(n5285), .B0(n544), .B1(n5306), .Y(n1511) );
  OAI22X1 U8076 ( .A0(n592), .A1(n5284), .B0(n640), .B1(n5306), .Y(n1644) );
  OAI22X1 U8077 ( .A0(n383), .A1(n5287), .B0(n431), .B1(n5305), .Y(n1241) );
  OAI22X1 U8078 ( .A0(n511), .A1(n5285), .B0(n543), .B1(n5306), .Y(n1507) );
  OAI22X1 U8079 ( .A0(n591), .A1(n5284), .B0(n639), .B1(n5307), .Y(n1640) );
  OAI22X1 U8080 ( .A0(n449), .A1(n5286), .B0(n481), .B1(n5305), .Y(n1383) );
  OAI22X1 U8081 ( .A0(n448), .A1(n5286), .B0(n480), .B1(n5305), .Y(n1379) );
  OAI22X1 U8082 ( .A0(n447), .A1(n5286), .B0(n479), .B1(n5305), .Y(n1375) );
  OAI22X1 U8083 ( .A0(n446), .A1(n5286), .B0(n478), .B1(n5305), .Y(n1371) );
  OAI22X1 U8084 ( .A0(n445), .A1(n5286), .B0(n477), .B1(n5304), .Y(n1367) );
  OAI22X1 U8085 ( .A0(n444), .A1(n5286), .B0(n476), .B1(n5305), .Y(n1363) );
  OAI22X1 U8086 ( .A0(n443), .A1(n5286), .B0(n475), .B1(n5305), .Y(n1359) );
  OAI22X1 U8087 ( .A0(n587), .A1(n5284), .B0(n635), .B1(n5307), .Y(n1624) );
  OAI22X1 U8088 ( .A0(n442), .A1(n5287), .B0(n474), .B1(n5305), .Y(n1355) );
  OAI22X1 U8089 ( .A0(n586), .A1(n5284), .B0(n634), .B1(n5306), .Y(n1620) );
  OAI22X1 U8090 ( .A0(n510), .A1(n5285), .B0(n542), .B1(n5306), .Y(n1503) );
  OAI22X1 U8091 ( .A0(n441), .A1(n5287), .B0(n473), .B1(n5305), .Y(n1351) );
  OAI22X1 U8092 ( .A0(n585), .A1(n5284), .B0(n633), .B1(n5307), .Y(n1616) );
  OAI22X1 U8093 ( .A0(n440), .A1(n5287), .B0(n472), .B1(n5305), .Y(n1347) );
  OAI22X1 U8094 ( .A0(n584), .A1(n5284), .B0(n632), .B1(n5307), .Y(n1612) );
  OAI22X1 U8095 ( .A0(n439), .A1(n5287), .B0(n471), .B1(n5305), .Y(n1343) );
  OAI22X1 U8096 ( .A0(n438), .A1(n5287), .B0(n470), .B1(n5305), .Y(n1339) );
  OAI22X1 U8097 ( .A0(n437), .A1(n5287), .B0(n469), .B1(n5305), .Y(n1335) );
  OAI22X1 U8098 ( .A0(n436), .A1(n5287), .B0(n468), .B1(n5305), .Y(n1331) );
  OAI22X1 U8099 ( .A0(n435), .A1(n5287), .B0(n467), .B1(n5305), .Y(n1327) );
  OAI22X1 U8100 ( .A0(n434), .A1(n5287), .B0(n466), .B1(n5305), .Y(n1323) );
  OAI22X1 U8101 ( .A0(n509), .A1(n5285), .B0(n541), .B1(n5306), .Y(n1499) );
  OAI22X1 U8102 ( .A0(n508), .A1(n5285), .B0(n540), .B1(n5306), .Y(n1495) );
  OAI22X1 U8103 ( .A0(n507), .A1(n5285), .B0(n539), .B1(n5306), .Y(n1491) );
  OAI22X1 U8104 ( .A0(n506), .A1(n5285), .B0(n538), .B1(n5306), .Y(n1487) );
  OAI22X1 U8105 ( .A0(n505), .A1(n5285), .B0(n537), .B1(n5306), .Y(n1483) );
  OAI22X1 U8106 ( .A0(n504), .A1(n5285), .B0(n536), .B1(n5307), .Y(n1479) );
  OAI22X1 U8107 ( .A0(n458), .A1(n5304), .B0(n490), .B1(n5264), .Y(n1289) );
  OAI22X1 U8108 ( .A0(n457), .A1(n5310), .B0(n489), .B1(n5264), .Y(n1285) );
  OAI22X1 U8109 ( .A0(n456), .A1(n5304), .B0(n488), .B1(n5264), .Y(n1281) );
  OAI22X1 U8110 ( .A0(n455), .A1(n5310), .B0(n487), .B1(n5264), .Y(n1277) );
  OAI22X1 U8111 ( .A0(n454), .A1(n5304), .B0(n486), .B1(n5264), .Y(n1273) );
  OAI22X1 U8112 ( .A0(n453), .A1(n5310), .B0(n485), .B1(n5264), .Y(n1269) );
  OAI22X1 U8113 ( .A0(n452), .A1(n5304), .B0(n484), .B1(n5264), .Y(n1265) );
  OAI22X1 U8114 ( .A0(n451), .A1(n5310), .B0(n483), .B1(n5264), .Y(n1261) );
  OAI22X1 U8115 ( .A0(n450), .A1(n5309), .B0(n482), .B1(n5264), .Y(n1256) );
  NOR2X1 U8116 ( .A(n1092), .B(store_cnt[0]), .Y(N14270) );
  NAND2X1 U8117 ( .A(c_plus[28]), .B(n824), .Y(n810) );
  AOI2BB1X1 U8118 ( .A0N(store_cnt[1]), .A1N(n1092), .B0(N14270), .Y(n1093) );
  NAND2X1 U8119 ( .A(c_plus[30]), .B(n837), .Y(n812) );
  NAND2X1 U8120 ( .A(c_plus[29]), .B(n837), .Y(n811) );
  OAI2BB1X1 U8121 ( .A0N(n1090), .A1N(store_cnt[3]), .B0(n1091), .Y(N14273) );
  OR4X2 U8122 ( .A(n866), .B(n1092), .C(n5896), .D(store_cnt[3]), .Y(n1091) );
  OAI21XL U8123 ( .A0(n1092), .A1(store_cnt[2]), .B0(n1093), .Y(n1090) );
  INVX1 U8124 ( .A(out_cnt[0]), .Y(n5971) );
  NOR3X1 U8125 ( .A(n5088), .B(n5087), .C(cal_cnt[0]), .Y(n1651) );
  NOR2X1 U8126 ( .A(n1007), .B(n1008), .Y(n1005) );
  XNOR2X1 U8127 ( .A(in_cnt[3]), .B(n5887), .Y(n1007) );
  XNOR2X1 U8128 ( .A(in_cnt[2]), .B(n5887), .Y(n1008) );
  BUFX3 U8129 ( .A(n1652), .Y(n5058) );
  NAND3X1 U8130 ( .A(n5087), .B(n5088), .C(cal_cnt[0]), .Y(n1652) );
  INVX1 U8131 ( .A(mem_weight_Q[16]), .Y(n5784) );
  INVX1 U8132 ( .A(mem_weight_Q[17]), .Y(n5783) );
  INVX1 U8133 ( .A(mem_weight_Q[18]), .Y(n5782) );
  INVX1 U8134 ( .A(mem_weight_Q[19]), .Y(n5781) );
  INVX1 U8135 ( .A(mem_weight_Q[20]), .Y(n5779) );
  INVX1 U8136 ( .A(mem_weight_Q[21]), .Y(n5778) );
  INVX1 U8137 ( .A(mem_weight_Q[22]), .Y(n5777) );
  INVX1 U8138 ( .A(mem_weight_Q[23]), .Y(n5776) );
  INVX1 U8139 ( .A(mem_weight_Q[24]), .Y(n5775) );
  INVX1 U8140 ( .A(mem_weight_Q[25]), .Y(n5774) );
  INVX1 U8141 ( .A(mem_weight_Q[26]), .Y(n5773) );
  INVX1 U8142 ( .A(mem_weight_Q[27]), .Y(n5772) );
  INVX1 U8143 ( .A(mem_weight_Q[28]), .Y(n5771) );
  INVX1 U8144 ( .A(mem_weight_Q[29]), .Y(n5770) );
  INVX1 U8145 ( .A(mem_weight_Q[30]), .Y(n5768) );
  INVX1 U8146 ( .A(mem_weight_Q[31]), .Y(n5767) );
  INVX1 U8147 ( .A(mem_weight_Q[0]), .Y(n5791) );
  INVX1 U8148 ( .A(mem_weight_Q[10]), .Y(n5790) );
  INVX1 U8149 ( .A(mem_weight_Q[11]), .Y(n5789) );
  INVX1 U8150 ( .A(mem_weight_Q[12]), .Y(n5788) );
  INVX1 U8151 ( .A(mem_weight_Q[13]), .Y(n5787) );
  INVX1 U8152 ( .A(mem_weight_Q[14]), .Y(n5786) );
  INVX1 U8153 ( .A(mem_weight_Q[15]), .Y(n5785) );
  INVX1 U8154 ( .A(mem_weight_Q[1]), .Y(n5780) );
  INVX1 U8155 ( .A(mem_weight_Q[2]), .Y(n5769) );
  INVX1 U8156 ( .A(mem_weight_Q[3]), .Y(n5758) );
  INVX1 U8157 ( .A(mem_weight_Q[4]), .Y(n5747) );
  INVX1 U8158 ( .A(mem_weight_Q[5]), .Y(n5736) );
  INVX1 U8159 ( .A(mem_weight_Q[6]), .Y(n5731) );
  INVX1 U8160 ( .A(mem_weight_Q[7]), .Y(n5730) );
  INVX1 U8161 ( .A(mem_weight_Q[8]), .Y(n5729) );
  INVX1 U8162 ( .A(mem_weight_Q[9]), .Y(n5728) );
  NAND2X1 U8163 ( .A(c_plus[27]), .B(n824), .Y(n809) );
  INVX1 U8164 ( .A(calin_cnt[2]), .Y(n5653) );
  INVX1 U8165 ( .A(mem_weight_Q[32]), .Y(n5766) );
  INVX1 U8166 ( .A(mem_weight_Q[33]), .Y(n5765) );
  INVX1 U8167 ( .A(mem_weight_Q[34]), .Y(n5764) );
  INVX1 U8168 ( .A(mem_weight_Q[35]), .Y(n5763) );
  INVX1 U8169 ( .A(mem_weight_Q[36]), .Y(n5762) );
  INVX1 U8170 ( .A(mem_weight_Q[37]), .Y(n5761) );
  INVX1 U8171 ( .A(mem_weight_Q[38]), .Y(n5760) );
  INVX1 U8172 ( .A(mem_weight_Q[39]), .Y(n5759) );
  INVX1 U8173 ( .A(mem_weight_Q[40]), .Y(n5757) );
  INVX1 U8174 ( .A(mem_weight_Q[41]), .Y(n5756) );
  INVX1 U8175 ( .A(mem_weight_Q[42]), .Y(n5755) );
  INVX1 U8176 ( .A(mem_weight_Q[43]), .Y(n5754) );
  INVX1 U8177 ( .A(mem_weight_Q[44]), .Y(n5753) );
  INVX1 U8178 ( .A(mem_weight_Q[45]), .Y(n5752) );
  INVX1 U8179 ( .A(mem_weight_Q[46]), .Y(n5751) );
  INVX1 U8180 ( .A(mem_weight_Q[47]), .Y(n5750) );
  INVX1 U8181 ( .A(mem_weight_Q[48]), .Y(n5749) );
  INVX1 U8182 ( .A(mem_weight_Q[49]), .Y(n5748) );
  INVX1 U8183 ( .A(mem_weight_Q[50]), .Y(n5746) );
  INVX1 U8184 ( .A(mem_weight_Q[51]), .Y(n5745) );
  INVX1 U8185 ( .A(mem_weight_Q[52]), .Y(n5744) );
  INVX1 U8186 ( .A(mem_weight_Q[53]), .Y(n5743) );
  INVX1 U8187 ( .A(mem_weight_Q[54]), .Y(n5742) );
  INVX1 U8188 ( .A(mem_weight_Q[55]), .Y(n5741) );
  INVX1 U8189 ( .A(mem_weight_Q[56]), .Y(n5740) );
  INVX1 U8190 ( .A(mem_weight_Q[57]), .Y(n5739) );
  INVX1 U8191 ( .A(mem_weight_Q[58]), .Y(n5738) );
  INVX1 U8192 ( .A(mem_weight_Q[59]), .Y(n5737) );
  INVX1 U8193 ( .A(mem_weight_Q[60]), .Y(n5735) );
  INVX1 U8194 ( .A(mem_weight_Q[61]), .Y(n5734) );
  INVX1 U8195 ( .A(mem_weight_Q[62]), .Y(n5733) );
  INVX1 U8196 ( .A(mem_weight_Q[63]), .Y(n5732) );
  INVX1 U8197 ( .A(mem_in_Q[0]), .Y(n5727) );
  INVX1 U8198 ( .A(mem_in_Q[10]), .Y(n5726) );
  INVX1 U8199 ( .A(mem_in_Q[11]), .Y(n5725) );
  INVX1 U8200 ( .A(mem_in_Q[12]), .Y(n5724) );
  INVX1 U8201 ( .A(mem_in_Q[13]), .Y(n5723) );
  INVX1 U8202 ( .A(mem_in_Q[14]), .Y(n5722) );
  INVX1 U8203 ( .A(mem_in_Q[15]), .Y(n5721) );
  INVX1 U8204 ( .A(mem_in_Q[1]), .Y(n5716) );
  INVX1 U8205 ( .A(mem_in_Q[2]), .Y(n5705) );
  INVX1 U8206 ( .A(mem_in_Q[3]), .Y(n5694) );
  INVX1 U8207 ( .A(mem_in_Q[4]), .Y(n5683) );
  INVX1 U8208 ( .A(mem_in_Q[5]), .Y(n5672) );
  INVX1 U8209 ( .A(mem_in_Q[6]), .Y(n5667) );
  INVX1 U8210 ( .A(mem_in_Q[7]), .Y(n5666) );
  INVX1 U8211 ( .A(mem_in_Q[8]), .Y(n5665) );
  INVX1 U8212 ( .A(mem_in_Q[9]), .Y(n5664) );
  INVX1 U8213 ( .A(mem_in_Q[48]), .Y(n5685) );
  INVX1 U8214 ( .A(mem_in_Q[49]), .Y(n5684) );
  INVX1 U8215 ( .A(mem_in_Q[50]), .Y(n5682) );
  INVX1 U8216 ( .A(mem_in_Q[51]), .Y(n5681) );
  INVX1 U8217 ( .A(mem_in_Q[52]), .Y(n5680) );
  INVX1 U8218 ( .A(mem_in_Q[53]), .Y(n5679) );
  INVX1 U8219 ( .A(mem_in_Q[54]), .Y(n5678) );
  INVX1 U8220 ( .A(mem_in_Q[55]), .Y(n5677) );
  INVX1 U8221 ( .A(mem_in_Q[56]), .Y(n5676) );
  INVX1 U8222 ( .A(mem_in_Q[57]), .Y(n5675) );
  INVX1 U8223 ( .A(mem_in_Q[58]), .Y(n5674) );
  INVX1 U8224 ( .A(mem_in_Q[59]), .Y(n5673) );
  INVX1 U8225 ( .A(mem_in_Q[60]), .Y(n5671) );
  INVX1 U8226 ( .A(mem_in_Q[61]), .Y(n5670) );
  INVX1 U8227 ( .A(mem_in_Q[62]), .Y(n5669) );
  INVX1 U8228 ( .A(mem_in_Q[63]), .Y(n5668) );
  INVX1 U8229 ( .A(mem_in_Q[32]), .Y(n5702) );
  INVX1 U8230 ( .A(mem_in_Q[33]), .Y(n5701) );
  INVX1 U8231 ( .A(mem_in_Q[34]), .Y(n5700) );
  INVX1 U8232 ( .A(mem_in_Q[35]), .Y(n5699) );
  INVX1 U8233 ( .A(mem_in_Q[36]), .Y(n5698) );
  INVX1 U8234 ( .A(mem_in_Q[37]), .Y(n5697) );
  INVX1 U8235 ( .A(mem_in_Q[38]), .Y(n5696) );
  INVX1 U8236 ( .A(mem_in_Q[39]), .Y(n5695) );
  INVX1 U8237 ( .A(mem_in_Q[40]), .Y(n5693) );
  INVX1 U8238 ( .A(mem_in_Q[41]), .Y(n5692) );
  INVX1 U8239 ( .A(mem_in_Q[42]), .Y(n5691) );
  INVX1 U8240 ( .A(mem_in_Q[43]), .Y(n5690) );
  INVX1 U8241 ( .A(mem_in_Q[44]), .Y(n5689) );
  INVX1 U8242 ( .A(mem_in_Q[45]), .Y(n5688) );
  INVX1 U8243 ( .A(mem_in_Q[46]), .Y(n5687) );
  INVX1 U8244 ( .A(mem_in_Q[47]), .Y(n5686) );
  XNOR2X1 U8245 ( .A(in_addr_cnt[8]), .B(N1234), .Y(n982) );
  INVX1 U8246 ( .A(n1035), .Y(n5837) );
  AOI22XL U8247 ( .A0(N14360), .A1(n1031), .B0(N14366), .B1(n1032), .Y(n1035)
         );
  OAI32X1 U8248 ( .A0(n1092), .A1(store_cnt[2]), .A2(n866), .B0(n1093), .B1(
        n5896), .Y(N14272) );
  BUFX3 U8249 ( .A(cal_cnt[1]), .Y(n5088) );
  AND2X2 U8250 ( .A(in_addr_cnt[0]), .B(n4495), .Y(n984) );
  XNOR2X1 U8251 ( .A(in_addr_cnt[6]), .B(N1232), .Y(n4495) );
  BUFX3 U8252 ( .A(cal_cnt[2]), .Y(n5087) );
  INVX1 U8253 ( .A(mem_in_Q[16]), .Y(n5720) );
  INVX1 U8254 ( .A(mem_in_Q[17]), .Y(n5719) );
  INVX1 U8255 ( .A(mem_in_Q[18]), .Y(n5718) );
  INVX1 U8256 ( .A(mem_in_Q[19]), .Y(n5717) );
  INVX1 U8257 ( .A(mem_in_Q[20]), .Y(n5715) );
  INVX1 U8258 ( .A(mem_in_Q[21]), .Y(n5714) );
  INVX1 U8259 ( .A(mem_in_Q[22]), .Y(n5713) );
  INVX1 U8260 ( .A(mem_in_Q[23]), .Y(n5712) );
  INVX1 U8261 ( .A(mem_in_Q[24]), .Y(n5711) );
  INVX1 U8262 ( .A(mem_in_Q[25]), .Y(n5710) );
  INVX1 U8263 ( .A(mem_in_Q[26]), .Y(n5709) );
  INVX1 U8264 ( .A(mem_in_Q[27]), .Y(n5708) );
  INVX1 U8265 ( .A(mem_in_Q[28]), .Y(n5707) );
  INVX1 U8266 ( .A(mem_in_Q[29]), .Y(n5706) );
  INVX1 U8267 ( .A(mem_in_Q[30]), .Y(n5704) );
  INVX1 U8268 ( .A(mem_in_Q[31]), .Y(n5703) );
  AOI31X1 U8269 ( .A0(n1206), .A1(n1207), .A2(n1208), .B0(n5316), .Y(N12070)
         );
  AOI22X1 U8270 ( .A0(n5060), .A1(x_matrix[10]), .B0(n1187), .B1(x_matrix[90]), 
        .Y(n1207) );
  AOI22X1 U8271 ( .A0(n5302), .A1(x_matrix[170]), .B0(n1189), .B1(
        x_matrix[266]), .Y(n1206) );
  AOI221X1 U8272 ( .A0(n5314), .A1(x_matrix[362]), .B0(n5270), .B1(
        x_matrix[458]), .C0(n1209), .Y(n1208) );
  AOI31X1 U8273 ( .A0(n1202), .A1(n1203), .A2(n1204), .B0(n5321), .Y(N12071)
         );
  AOI22X1 U8274 ( .A0(n5060), .A1(x_matrix[11]), .B0(n1187), .B1(x_matrix[91]), 
        .Y(n1203) );
  AOI22X1 U8275 ( .A0(n5302), .A1(x_matrix[171]), .B0(n1189), .B1(
        x_matrix[267]), .Y(n1202) );
  AOI221X1 U8276 ( .A0(n5314), .A1(x_matrix[363]), .B0(n5266), .B1(
        x_matrix[459]), .C0(n1205), .Y(n1204) );
  AOI31X1 U8277 ( .A0(n1198), .A1(n1199), .A2(n1200), .B0(n5316), .Y(N12072)
         );
  AOI22X1 U8278 ( .A0(n5060), .A1(x_matrix[12]), .B0(n1187), .B1(x_matrix[92]), 
        .Y(n1199) );
  AOI22X1 U8279 ( .A0(n5302), .A1(x_matrix[172]), .B0(n1189), .B1(
        x_matrix[268]), .Y(n1198) );
  AOI221X1 U8280 ( .A0(n5314), .A1(x_matrix[364]), .B0(n5269), .B1(
        x_matrix[460]), .C0(n1201), .Y(n1200) );
  AOI31X1 U8281 ( .A0(n1194), .A1(n1195), .A2(n1196), .B0(n5321), .Y(N12073)
         );
  AOI22X1 U8282 ( .A0(n5060), .A1(x_matrix[13]), .B0(n1187), .B1(x_matrix[93]), 
        .Y(n1195) );
  AOI22X1 U8283 ( .A0(n1188), .A1(x_matrix[173]), .B0(n1189), .B1(
        x_matrix[269]), .Y(n1194) );
  AOI221X1 U8284 ( .A0(n5314), .A1(x_matrix[365]), .B0(n5266), .B1(
        x_matrix[461]), .C0(n1197), .Y(n1196) );
  AOI31X1 U8285 ( .A0(n1190), .A1(n1191), .A2(n1192), .B0(n5316), .Y(N12074)
         );
  AOI22X1 U8286 ( .A0(n5060), .A1(x_matrix[14]), .B0(n1187), .B1(x_matrix[94]), 
        .Y(n1191) );
  AOI22X1 U8287 ( .A0(n1188), .A1(x_matrix[174]), .B0(n1189), .B1(
        x_matrix[270]), .Y(n1190) );
  AOI221X1 U8288 ( .A0(n5314), .A1(x_matrix[366]), .B0(n5272), .B1(
        x_matrix[462]), .C0(n1193), .Y(n1192) );
  AOI31X1 U8289 ( .A0(n1179), .A1(n1180), .A2(n1181), .B0(n5321), .Y(N12075)
         );
  AOI22X1 U8290 ( .A0(n5060), .A1(x_matrix[15]), .B0(n1187), .B1(x_matrix[95]), 
        .Y(n1180) );
  AOI22X1 U8291 ( .A0(n5302), .A1(x_matrix[175]), .B0(n1189), .B1(
        x_matrix[271]), .Y(n1179) );
  AOI221X1 U8292 ( .A0(n5314), .A1(x_matrix[367]), .B0(n5275), .B1(
        x_matrix[463]), .C0(n1184), .Y(n1181) );
  AOI31X1 U8293 ( .A0(n1214), .A1(n1215), .A2(n1216), .B0(n5316), .Y(N12068)
         );
  AOI22X1 U8294 ( .A0(n5060), .A1(x_matrix[8]), .B0(n1187), .B1(x_matrix[88]), 
        .Y(n1215) );
  AOI22X1 U8295 ( .A0(n1188), .A1(x_matrix[168]), .B0(n1189), .B1(
        x_matrix[264]), .Y(n1214) );
  AOI221X1 U8296 ( .A0(n5314), .A1(x_matrix[360]), .B0(n5271), .B1(
        x_matrix[456]), .C0(n1217), .Y(n1216) );
  AOI31X1 U8297 ( .A0(n1210), .A1(n1211), .A2(n1212), .B0(n5321), .Y(N12069)
         );
  AOI22X1 U8298 ( .A0(n5060), .A1(x_matrix[9]), .B0(n1187), .B1(x_matrix[89]), 
        .Y(n1211) );
  AOI22X1 U8299 ( .A0(n1188), .A1(x_matrix[169]), .B0(n1189), .B1(
        x_matrix[265]), .Y(n1210) );
  AOI221X1 U8300 ( .A0(n5314), .A1(x_matrix[361]), .B0(n5267), .B1(
        x_matrix[457]), .C0(n1213), .Y(n1212) );
  AOI31X1 U8301 ( .A0(n1645), .A1(n1646), .A2(n1647), .B0(n5316), .Y(N11490)
         );
  AOI22X1 U8302 ( .A0(n1522), .A1(x_matrix[624]), .B0(n5059), .B1(
        x_matrix[736]), .Y(n1645) );
  AOI22X1 U8303 ( .A0(n5253), .A1(x_matrix[416]), .B0(n1455), .B1(
        x_matrix[512]), .Y(n1646) );
  AOI221X1 U8304 ( .A0(n5282), .A1(x_matrix[224]), .B0(n1322), .B1(
        x_matrix[320]), .C0(n1650), .Y(n1647) );
  AOI31X1 U8305 ( .A0(n1605), .A1(n1606), .A2(n1607), .B0(n5316), .Y(N11500)
         );
  AOI22X1 U8306 ( .A0(n1522), .A1(x_matrix[634]), .B0(n5059), .B1(
        x_matrix[746]), .Y(n1605) );
  AOI22X1 U8307 ( .A0(n5253), .A1(x_matrix[426]), .B0(n5251), .B1(
        x_matrix[522]), .Y(n1606) );
  AOI221X1 U8308 ( .A0(n5282), .A1(x_matrix[234]), .B0(n5259), .B1(
        x_matrix[330]), .C0(n1608), .Y(n1607) );
  AOI31X1 U8309 ( .A0(n1601), .A1(n1602), .A2(n1603), .B0(n5316), .Y(N11501)
         );
  AOI22X1 U8310 ( .A0(n1522), .A1(x_matrix[635]), .B0(n5059), .B1(
        x_matrix[747]), .Y(n1601) );
  AOI22X1 U8311 ( .A0(n5253), .A1(x_matrix[427]), .B0(n1455), .B1(
        x_matrix[523]), .Y(n1602) );
  AOI221X1 U8312 ( .A0(n5282), .A1(x_matrix[235]), .B0(n5259), .B1(
        x_matrix[331]), .C0(n1604), .Y(n1603) );
  AOI31X1 U8313 ( .A0(n1597), .A1(n1598), .A2(n1599), .B0(n5316), .Y(N11502)
         );
  AOI22X1 U8314 ( .A0(n1522), .A1(x_matrix[636]), .B0(n5059), .B1(
        x_matrix[748]), .Y(n1597) );
  AOI22X1 U8315 ( .A0(n5254), .A1(x_matrix[428]), .B0(n1455), .B1(
        x_matrix[524]), .Y(n1598) );
  AOI221X1 U8316 ( .A0(n5282), .A1(x_matrix[236]), .B0(n5259), .B1(
        x_matrix[332]), .C0(n1600), .Y(n1599) );
  AOI31X1 U8317 ( .A0(n1641), .A1(n1642), .A2(n1643), .B0(n5316), .Y(N11491)
         );
  AOI22X1 U8318 ( .A0(n1522), .A1(x_matrix[625]), .B0(n5059), .B1(
        x_matrix[737]), .Y(n1641) );
  AOI22X1 U8319 ( .A0(n5253), .A1(x_matrix[417]), .B0(n5251), .B1(
        x_matrix[513]), .Y(n1642) );
  AOI221X1 U8320 ( .A0(n5282), .A1(x_matrix[225]), .B0(n5259), .B1(
        x_matrix[321]), .C0(n1644), .Y(n1643) );
  AOI31X1 U8321 ( .A0(n1637), .A1(n1638), .A2(n1639), .B0(n5316), .Y(N11492)
         );
  AOI22X1 U8322 ( .A0(n1522), .A1(x_matrix[626]), .B0(n5059), .B1(
        x_matrix[738]), .Y(n1637) );
  AOI22X1 U8323 ( .A0(n5254), .A1(x_matrix[418]), .B0(n5251), .B1(
        x_matrix[514]), .Y(n1638) );
  AOI221X1 U8324 ( .A0(n5282), .A1(x_matrix[226]), .B0(n5259), .B1(
        x_matrix[322]), .C0(n1640), .Y(n1639) );
  AOI31X1 U8325 ( .A0(n1633), .A1(n1634), .A2(n1635), .B0(n5316), .Y(N11493)
         );
  AOI22X1 U8326 ( .A0(n1522), .A1(x_matrix[627]), .B0(n5059), .B1(
        x_matrix[739]), .Y(n1633) );
  AOI22X1 U8327 ( .A0(n1389), .A1(x_matrix[419]), .B0(n5251), .B1(
        x_matrix[515]), .Y(n1634) );
  AOI221X1 U8328 ( .A0(n5282), .A1(x_matrix[227]), .B0(n5259), .B1(
        x_matrix[323]), .C0(n1636), .Y(n1635) );
  AOI31X1 U8329 ( .A0(n1629), .A1(n1630), .A2(n1631), .B0(n5316), .Y(N11494)
         );
  AOI22X1 U8330 ( .A0(n1522), .A1(x_matrix[628]), .B0(n5059), .B1(
        x_matrix[740]), .Y(n1629) );
  AOI22X1 U8331 ( .A0(n1389), .A1(x_matrix[420]), .B0(n5251), .B1(
        x_matrix[516]), .Y(n1630) );
  AOI221X1 U8332 ( .A0(n5282), .A1(x_matrix[228]), .B0(n5259), .B1(
        x_matrix[324]), .C0(n1632), .Y(n1631) );
  AOI31X1 U8333 ( .A0(n1625), .A1(n1626), .A2(n1627), .B0(n5316), .Y(N11495)
         );
  AOI22X1 U8334 ( .A0(n1522), .A1(x_matrix[629]), .B0(n5059), .B1(
        x_matrix[741]), .Y(n1625) );
  AOI22X1 U8335 ( .A0(n5254), .A1(x_matrix[421]), .B0(n5251), .B1(
        x_matrix[517]), .Y(n1626) );
  AOI221X1 U8336 ( .A0(n5282), .A1(x_matrix[229]), .B0(n5259), .B1(
        x_matrix[325]), .C0(n1628), .Y(n1627) );
  AOI31X1 U8337 ( .A0(n1621), .A1(n1622), .A2(n1623), .B0(n5316), .Y(N11496)
         );
  AOI22X1 U8338 ( .A0(n1522), .A1(x_matrix[630]), .B0(n5059), .B1(
        x_matrix[742]), .Y(n1621) );
  AOI22X1 U8339 ( .A0(n1389), .A1(x_matrix[422]), .B0(n5251), .B1(
        x_matrix[518]), .Y(n1622) );
  AOI221X1 U8340 ( .A0(n5282), .A1(x_matrix[230]), .B0(n5259), .B1(
        x_matrix[326]), .C0(n1624), .Y(n1623) );
  AOI31X1 U8341 ( .A0(n1617), .A1(n1618), .A2(n1619), .B0(n5316), .Y(N11497)
         );
  AOI22X1 U8342 ( .A0(n1522), .A1(x_matrix[631]), .B0(n5059), .B1(
        x_matrix[743]), .Y(n1617) );
  AOI22X1 U8343 ( .A0(n1389), .A1(x_matrix[423]), .B0(n5251), .B1(
        x_matrix[519]), .Y(n1618) );
  AOI221X1 U8344 ( .A0(n5282), .A1(x_matrix[231]), .B0(n5259), .B1(
        x_matrix[327]), .C0(n1620), .Y(n1619) );
  AOI31X1 U8345 ( .A0(n1613), .A1(n1614), .A2(n1615), .B0(n5316), .Y(N11498)
         );
  AOI22X1 U8346 ( .A0(n1522), .A1(x_matrix[632]), .B0(n5059), .B1(
        x_matrix[744]), .Y(n1613) );
  AOI22X1 U8347 ( .A0(n1389), .A1(x_matrix[424]), .B0(n5251), .B1(
        x_matrix[520]), .Y(n1614) );
  AOI221X1 U8348 ( .A0(n5282), .A1(x_matrix[232]), .B0(n5259), .B1(
        x_matrix[328]), .C0(n1616), .Y(n1615) );
  AOI31X1 U8349 ( .A0(n1609), .A1(n1610), .A2(n1611), .B0(n5316), .Y(N11499)
         );
  AOI22X1 U8350 ( .A0(n1522), .A1(x_matrix[633]), .B0(n5059), .B1(
        x_matrix[745]), .Y(n1609) );
  AOI22X1 U8351 ( .A0(n1389), .A1(x_matrix[425]), .B0(n5251), .B1(
        x_matrix[521]), .Y(n1610) );
  AOI221X1 U8352 ( .A0(n5282), .A1(x_matrix[233]), .B0(n5259), .B1(
        x_matrix[329]), .C0(n1612), .Y(n1611) );
  AOI31X1 U8353 ( .A0(n1246), .A1(n1247), .A2(n1248), .B0(n5321), .Y(N12060)
         );
  AOI22X1 U8354 ( .A0(n5060), .A1(x_matrix[0]), .B0(n1187), .B1(x_matrix[80]), 
        .Y(n1247) );
  AOI22X1 U8355 ( .A0(n5302), .A1(x_matrix[160]), .B0(n5298), .B1(
        x_matrix[256]), .Y(n1246) );
  AOI221X1 U8356 ( .A0(n5314), .A1(x_matrix[352]), .B0(n5271), .B1(
        x_matrix[448]), .C0(n1249), .Y(n1248) );
  AOI31X1 U8357 ( .A0(n1512), .A1(n1513), .A2(n1514), .B0(n5318), .Y(N11681)
         );
  AOI22X1 U8358 ( .A0(n5253), .A1(x_matrix[592]), .B0(n1455), .B1(
        x_matrix[704]), .Y(n1512) );
  AOI22X1 U8359 ( .A0(n5282), .A1(x_matrix[384]), .B0(n5258), .B1(
        x_matrix[480]), .Y(n1513) );
  AOI221X1 U8360 ( .A0(n5314), .A1(x_matrix[64]), .B0(n5265), .B1(
        x_matrix[144]), .C0(n1515), .Y(n1514) );
  AOI31X1 U8361 ( .A0(n1472), .A1(n1473), .A2(n1474), .B0(n5317), .Y(N11691)
         );
  AOI22X1 U8362 ( .A0(n1389), .A1(x_matrix[602]), .B0(n1455), .B1(
        x_matrix[714]), .Y(n1472) );
  AOI22X1 U8363 ( .A0(n5282), .A1(x_matrix[394]), .B0(n1322), .B1(
        x_matrix[490]), .Y(n1473) );
  AOI221X1 U8364 ( .A0(n5314), .A1(x_matrix[74]), .B0(n5276), .B1(
        x_matrix[154]), .C0(n1475), .Y(n1474) );
  AOI31X1 U8365 ( .A0(n1468), .A1(n1469), .A2(n1470), .B0(n5318), .Y(N11692)
         );
  AOI22X1 U8366 ( .A0(n5253), .A1(x_matrix[603]), .B0(n1455), .B1(
        x_matrix[715]), .Y(n1468) );
  AOI22X1 U8367 ( .A0(n5282), .A1(x_matrix[395]), .B0(n1322), .B1(
        x_matrix[491]), .Y(n1469) );
  AOI221X1 U8368 ( .A0(n5314), .A1(x_matrix[75]), .B0(n5275), .B1(
        x_matrix[155]), .C0(n1471), .Y(n1470) );
  AOI31X1 U8369 ( .A0(n1464), .A1(n1465), .A2(n1466), .B0(n5317), .Y(N11693)
         );
  AOI22X1 U8370 ( .A0(n1389), .A1(x_matrix[604]), .B0(n1455), .B1(
        x_matrix[716]), .Y(n1464) );
  AOI22X1 U8371 ( .A0(n5282), .A1(x_matrix[396]), .B0(n1322), .B1(
        x_matrix[492]), .Y(n1465) );
  AOI221X1 U8372 ( .A0(n5314), .A1(x_matrix[76]), .B0(n5275), .B1(
        x_matrix[156]), .C0(n1467), .Y(n1466) );
  AOI31X1 U8373 ( .A0(n1460), .A1(n1461), .A2(n1462), .B0(n5318), .Y(N11694)
         );
  AOI22X1 U8374 ( .A0(n1389), .A1(x_matrix[605]), .B0(n1455), .B1(
        x_matrix[717]), .Y(n1460) );
  AOI22X1 U8375 ( .A0(n5282), .A1(x_matrix[397]), .B0(n1322), .B1(
        x_matrix[493]), .Y(n1461) );
  AOI221X1 U8376 ( .A0(n5314), .A1(x_matrix[77]), .B0(n5275), .B1(
        x_matrix[157]), .C0(n1463), .Y(n1462) );
  AOI31X1 U8377 ( .A0(n1593), .A1(n1594), .A2(n1595), .B0(n5317), .Y(N11503)
         );
  AOI22X1 U8378 ( .A0(n1522), .A1(x_matrix[637]), .B0(n5059), .B1(
        x_matrix[749]), .Y(n1593) );
  AOI22X1 U8379 ( .A0(n5253), .A1(x_matrix[429]), .B0(n1455), .B1(
        x_matrix[525]), .Y(n1594) );
  AOI221X1 U8380 ( .A0(n5282), .A1(x_matrix[237]), .B0(n5259), .B1(
        x_matrix[333]), .C0(n1596), .Y(n1595) );
  AOI31X1 U8381 ( .A0(n1456), .A1(n1457), .A2(n1458), .B0(n5317), .Y(N11695)
         );
  AOI22X1 U8382 ( .A0(n1389), .A1(x_matrix[606]), .B0(n1455), .B1(
        x_matrix[718]), .Y(n1456) );
  AOI22X1 U8383 ( .A0(n5282), .A1(x_matrix[398]), .B0(n1322), .B1(
        x_matrix[494]), .Y(n1457) );
  AOI221X1 U8384 ( .A0(n5314), .A1(x_matrix[78]), .B0(n5275), .B1(
        x_matrix[158]), .C0(n1459), .Y(n1458) );
  AOI31X1 U8385 ( .A0(n1589), .A1(n1590), .A2(n1591), .B0(n5317), .Y(N11504)
         );
  AOI22X1 U8386 ( .A0(n1522), .A1(x_matrix[638]), .B0(n5059), .B1(
        x_matrix[750]), .Y(n1589) );
  AOI22X1 U8387 ( .A0(n5253), .A1(x_matrix[430]), .B0(n1455), .B1(
        x_matrix[526]), .Y(n1590) );
  AOI221X1 U8388 ( .A0(n5282), .A1(x_matrix[238]), .B0(n5259), .B1(
        x_matrix[334]), .C0(n1592), .Y(n1591) );
  AOI31X1 U8389 ( .A0(n1451), .A1(n1452), .A2(n1453), .B0(n5318), .Y(N11696)
         );
  AOI22X1 U8390 ( .A0(n5253), .A1(x_matrix[607]), .B0(n1455), .B1(
        x_matrix[719]), .Y(n1451) );
  AOI22X1 U8391 ( .A0(n5282), .A1(x_matrix[399]), .B0(n1322), .B1(
        x_matrix[495]), .Y(n1452) );
  AOI221X1 U8392 ( .A0(n1183), .A1(x_matrix[79]), .B0(n5275), .B1(
        x_matrix[159]), .C0(n1454), .Y(n1453) );
  AOI31X1 U8393 ( .A0(n1584), .A1(n1585), .A2(n1586), .B0(n5317), .Y(N11505)
         );
  AOI22X1 U8394 ( .A0(n1522), .A1(x_matrix[639]), .B0(n5059), .B1(
        x_matrix[751]), .Y(n1584) );
  AOI22X1 U8395 ( .A0(n5253), .A1(x_matrix[431]), .B0(n1455), .B1(
        x_matrix[527]), .Y(n1585) );
  AOI221X1 U8396 ( .A0(n5282), .A1(x_matrix[239]), .B0(n5259), .B1(
        x_matrix[335]), .C0(n1587), .Y(n1586) );
  AOI31X1 U8397 ( .A0(n1314), .A1(n1315), .A2(n1316), .B0(n5320), .Y(N11964)
         );
  AOI22X1 U8398 ( .A0(n1187), .A1(x_matrix[16]), .B0(n1188), .B1(x_matrix[96]), 
        .Y(n1315) );
  AOI22X1 U8399 ( .A0(n5298), .A1(x_matrix[176]), .B0(n5314), .B1(
        x_matrix[272]), .Y(n1314) );
  AOI221X1 U8400 ( .A0(n5293), .A1(x_matrix[544]), .B0(n1255), .B1(
        x_matrix[656]), .C0(n1317), .Y(n1316) );
  AOI31X1 U8401 ( .A0(n1579), .A1(n1580), .A2(n1581), .B0(n5317), .Y(N11584)
         );
  AOI22X1 U8402 ( .A0(n5251), .A1(x_matrix[608]), .B0(n1522), .B1(
        x_matrix[720]), .Y(n1579) );
  AOI22X1 U8403 ( .A0(n5257), .A1(x_matrix[400]), .B0(n5254), .B1(
        x_matrix[496]), .Y(n1580) );
  AOI221X1 U8404 ( .A0(n5289), .A1(x_matrix[208]), .B0(n1255), .B1(
        x_matrix[304]), .C0(n1582), .Y(n1581) );
  AOI31X1 U8405 ( .A0(n1310), .A1(n1311), .A2(n1312), .B0(n5320), .Y(N11965)
         );
  AOI22X1 U8406 ( .A0(n1187), .A1(x_matrix[17]), .B0(n1188), .B1(x_matrix[97]), 
        .Y(n1311) );
  AOI22X1 U8407 ( .A0(n1189), .A1(x_matrix[177]), .B0(n1183), .B1(
        x_matrix[273]), .Y(n1310) );
  AOI221X1 U8408 ( .A0(n5291), .A1(x_matrix[545]), .B0(n1255), .B1(
        x_matrix[657]), .C0(n1313), .Y(n1312) );
  AOI31X1 U8409 ( .A0(n1575), .A1(n1576), .A2(n1577), .B0(n5317), .Y(N11585)
         );
  AOI22X1 U8410 ( .A0(n5251), .A1(x_matrix[609]), .B0(n1522), .B1(
        x_matrix[721]), .Y(n1575) );
  AOI22X1 U8411 ( .A0(n5257), .A1(x_matrix[401]), .B0(n5254), .B1(
        x_matrix[497]), .Y(n1576) );
  AOI221X1 U8412 ( .A0(n5294), .A1(x_matrix[209]), .B0(n5282), .B1(
        x_matrix[305]), .C0(n1578), .Y(n1577) );
  AOI31X1 U8413 ( .A0(n1306), .A1(n1307), .A2(n1308), .B0(n5320), .Y(N11966)
         );
  AOI22X1 U8414 ( .A0(n1187), .A1(x_matrix[18]), .B0(n1188), .B1(x_matrix[98]), 
        .Y(n1307) );
  AOI22X1 U8415 ( .A0(n5298), .A1(x_matrix[178]), .B0(n5314), .B1(
        x_matrix[274]), .Y(n1306) );
  AOI221X1 U8416 ( .A0(n5292), .A1(x_matrix[546]), .B0(n5282), .B1(
        x_matrix[658]), .C0(n1309), .Y(n1308) );
  AOI31X1 U8417 ( .A0(n1571), .A1(n1572), .A2(n1573), .B0(n5317), .Y(N11586)
         );
  AOI22X1 U8418 ( .A0(n1455), .A1(x_matrix[610]), .B0(n1522), .B1(
        x_matrix[722]), .Y(n1571) );
  AOI22X1 U8419 ( .A0(n5257), .A1(x_matrix[402]), .B0(n5254), .B1(
        x_matrix[498]), .Y(n1572) );
  AOI221X1 U8420 ( .A0(n5296), .A1(x_matrix[210]), .B0(n5282), .B1(
        x_matrix[306]), .C0(n1574), .Y(n1573) );
  AOI31X1 U8421 ( .A0(n1302), .A1(n1303), .A2(n1304), .B0(n5320), .Y(N11967)
         );
  AOI22X1 U8422 ( .A0(n1187), .A1(x_matrix[19]), .B0(n1188), .B1(x_matrix[99]), 
        .Y(n1303) );
  AOI22X1 U8423 ( .A0(n1189), .A1(x_matrix[179]), .B0(n1183), .B1(
        x_matrix[275]), .Y(n1302) );
  AOI221X1 U8424 ( .A0(n5292), .A1(x_matrix[547]), .B0(n5282), .B1(
        x_matrix[659]), .C0(n1305), .Y(n1304) );
  AOI31X1 U8425 ( .A0(n1567), .A1(n1568), .A2(n1569), .B0(n5317), .Y(N11587)
         );
  AOI22X1 U8426 ( .A0(n5251), .A1(x_matrix[611]), .B0(n1522), .B1(
        x_matrix[723]), .Y(n1567) );
  AOI22X1 U8427 ( .A0(n5257), .A1(x_matrix[403]), .B0(n5254), .B1(
        x_matrix[499]), .Y(n1568) );
  AOI221X1 U8428 ( .A0(n5290), .A1(x_matrix[211]), .B0(n5282), .B1(
        x_matrix[307]), .C0(n1570), .Y(n1569) );
  AOI31X1 U8429 ( .A0(n1242), .A1(n1243), .A2(n1244), .B0(n5321), .Y(N12061)
         );
  AOI22X1 U8430 ( .A0(n5060), .A1(x_matrix[1]), .B0(n1187), .B1(x_matrix[81]), 
        .Y(n1243) );
  AOI22X1 U8431 ( .A0(n5302), .A1(x_matrix[161]), .B0(n1189), .B1(
        x_matrix[257]), .Y(n1242) );
  AOI221X1 U8432 ( .A0(n5314), .A1(x_matrix[353]), .B0(n5267), .B1(
        x_matrix[449]), .C0(n1245), .Y(n1244) );
  AOI31X1 U8433 ( .A0(n1508), .A1(n1509), .A2(n1510), .B0(n5318), .Y(N11682)
         );
  AOI22X1 U8434 ( .A0(n5253), .A1(x_matrix[593]), .B0(n1455), .B1(
        x_matrix[705]), .Y(n1508) );
  AOI22X1 U8435 ( .A0(n5282), .A1(x_matrix[385]), .B0(n5258), .B1(
        x_matrix[481]), .Y(n1509) );
  AOI221X1 U8436 ( .A0(n1183), .A1(x_matrix[65]), .B0(n5277), .B1(
        x_matrix[145]), .C0(n1511), .Y(n1510) );
  AOI31X1 U8437 ( .A0(n1298), .A1(n1299), .A2(n1300), .B0(n5320), .Y(N11968)
         );
  AOI22X1 U8438 ( .A0(n1187), .A1(x_matrix[20]), .B0(n1188), .B1(x_matrix[100]), .Y(n1299) );
  AOI22X1 U8439 ( .A0(n5298), .A1(x_matrix[180]), .B0(n5314), .B1(
        x_matrix[276]), .Y(n1298) );
  AOI221X1 U8440 ( .A0(n5291), .A1(x_matrix[548]), .B0(n5282), .B1(
        x_matrix[660]), .C0(n1301), .Y(n1300) );
  AOI31X1 U8441 ( .A0(n1563), .A1(n1564), .A2(n1565), .B0(n5317), .Y(N11588)
         );
  AOI22X1 U8442 ( .A0(n1455), .A1(x_matrix[612]), .B0(n1522), .B1(
        x_matrix[724]), .Y(n1563) );
  AOI22X1 U8443 ( .A0(n5258), .A1(x_matrix[404]), .B0(n5254), .B1(
        x_matrix[500]), .Y(n1564) );
  AOI221X1 U8444 ( .A0(n5296), .A1(x_matrix[212]), .B0(n5282), .B1(
        x_matrix[308]), .C0(n1566), .Y(n1565) );
  AOI31X1 U8445 ( .A0(n1294), .A1(n1295), .A2(n1296), .B0(n5320), .Y(N11969)
         );
  AOI22X1 U8446 ( .A0(n1187), .A1(x_matrix[21]), .B0(n1188), .B1(x_matrix[101]), .Y(n1295) );
  AOI22X1 U8447 ( .A0(n5298), .A1(x_matrix[181]), .B0(n1183), .B1(
        x_matrix[277]), .Y(n1294) );
  AOI221X1 U8448 ( .A0(n5292), .A1(x_matrix[549]), .B0(n5282), .B1(
        x_matrix[661]), .C0(n1297), .Y(n1296) );
  AOI31X1 U8449 ( .A0(n1559), .A1(n1560), .A2(n1561), .B0(n5317), .Y(N11589)
         );
  AOI22X1 U8450 ( .A0(n5251), .A1(x_matrix[613]), .B0(n1522), .B1(
        x_matrix[725]), .Y(n1559) );
  AOI22X1 U8451 ( .A0(n5257), .A1(x_matrix[405]), .B0(n5254), .B1(
        x_matrix[501]), .Y(n1560) );
  AOI221X1 U8452 ( .A0(n5288), .A1(x_matrix[213]), .B0(n5282), .B1(
        x_matrix[309]), .C0(n1562), .Y(n1561) );
  AOI31X1 U8453 ( .A0(n1290), .A1(n1291), .A2(n1292), .B0(n5320), .Y(N11970)
         );
  AOI22X1 U8454 ( .A0(n1187), .A1(x_matrix[22]), .B0(n1188), .B1(x_matrix[102]), .Y(n1291) );
  AOI22X1 U8455 ( .A0(n5298), .A1(x_matrix[182]), .B0(n5314), .B1(
        x_matrix[278]), .Y(n1290) );
  AOI221X1 U8456 ( .A0(n5290), .A1(x_matrix[550]), .B0(n5282), .B1(
        x_matrix[662]), .C0(n1293), .Y(n1292) );
  AOI31X1 U8457 ( .A0(n1555), .A1(n1556), .A2(n1557), .B0(n5317), .Y(N11590)
         );
  AOI22X1 U8458 ( .A0(n1455), .A1(x_matrix[614]), .B0(n1522), .B1(
        x_matrix[726]), .Y(n1555) );
  AOI22X1 U8459 ( .A0(n5258), .A1(x_matrix[406]), .B0(n5254), .B1(
        x_matrix[502]), .Y(n1556) );
  AOI221X1 U8460 ( .A0(n5296), .A1(x_matrix[214]), .B0(n5282), .B1(
        x_matrix[310]), .C0(n1558), .Y(n1557) );
  AOI31X1 U8461 ( .A0(n1286), .A1(n1287), .A2(n1288), .B0(n5320), .Y(N11971)
         );
  AOI22X1 U8462 ( .A0(n1187), .A1(x_matrix[23]), .B0(n1188), .B1(x_matrix[103]), .Y(n1287) );
  AOI22X1 U8463 ( .A0(n1189), .A1(x_matrix[183]), .B0(n1183), .B1(
        x_matrix[279]), .Y(n1286) );
  AOI221X1 U8464 ( .A0(n5290), .A1(x_matrix[551]), .B0(n5282), .B1(
        x_matrix[663]), .C0(n1289), .Y(n1288) );
  AOI31X1 U8465 ( .A0(n1551), .A1(n1552), .A2(n1553), .B0(n5317), .Y(N11591)
         );
  AOI22X1 U8466 ( .A0(n5251), .A1(x_matrix[615]), .B0(n1522), .B1(
        x_matrix[727]), .Y(n1551) );
  AOI22X1 U8467 ( .A0(n5257), .A1(x_matrix[407]), .B0(n5254), .B1(
        x_matrix[503]), .Y(n1552) );
  AOI221X1 U8468 ( .A0(n5296), .A1(x_matrix[215]), .B0(n5282), .B1(
        x_matrix[311]), .C0(n1554), .Y(n1553) );
  AOI31X1 U8469 ( .A0(n1282), .A1(n1283), .A2(n1284), .B0(n5320), .Y(N11972)
         );
  AOI22X1 U8470 ( .A0(n1187), .A1(x_matrix[24]), .B0(n1188), .B1(x_matrix[104]), .Y(n1283) );
  AOI22X1 U8471 ( .A0(n5298), .A1(x_matrix[184]), .B0(n5314), .B1(
        x_matrix[280]), .Y(n1282) );
  AOI221X1 U8472 ( .A0(n5292), .A1(x_matrix[552]), .B0(n5282), .B1(
        x_matrix[664]), .C0(n1285), .Y(n1284) );
  AOI31X1 U8473 ( .A0(n1547), .A1(n1548), .A2(n1549), .B0(n5317), .Y(N11592)
         );
  AOI22X1 U8474 ( .A0(n1455), .A1(x_matrix[616]), .B0(n1522), .B1(
        x_matrix[728]), .Y(n1547) );
  AOI22X1 U8475 ( .A0(n5258), .A1(x_matrix[408]), .B0(n5254), .B1(
        x_matrix[504]), .Y(n1548) );
  AOI221X1 U8476 ( .A0(n5296), .A1(x_matrix[216]), .B0(n5282), .B1(
        x_matrix[312]), .C0(n1550), .Y(n1549) );
  AOI31X1 U8477 ( .A0(n1278), .A1(n1279), .A2(n1280), .B0(n5320), .Y(N11973)
         );
  AOI22X1 U8478 ( .A0(n1187), .A1(x_matrix[25]), .B0(n1188), .B1(x_matrix[105]), .Y(n1279) );
  AOI22X1 U8479 ( .A0(n5298), .A1(x_matrix[185]), .B0(n1183), .B1(
        x_matrix[281]), .Y(n1278) );
  AOI221X1 U8480 ( .A0(n5290), .A1(x_matrix[553]), .B0(n5282), .B1(
        x_matrix[665]), .C0(n1281), .Y(n1280) );
  AOI31X1 U8481 ( .A0(n1543), .A1(n1544), .A2(n1545), .B0(n5317), .Y(N11593)
         );
  AOI22X1 U8482 ( .A0(n5251), .A1(x_matrix[617]), .B0(n1522), .B1(
        x_matrix[729]), .Y(n1543) );
  AOI22X1 U8483 ( .A0(n5257), .A1(x_matrix[409]), .B0(n5254), .B1(
        x_matrix[505]), .Y(n1544) );
  AOI221X1 U8484 ( .A0(n5295), .A1(x_matrix[217]), .B0(n5282), .B1(
        x_matrix[313]), .C0(n1546), .Y(n1545) );
  AOI31X1 U8485 ( .A0(n1274), .A1(n1275), .A2(n1276), .B0(n5320), .Y(N11974)
         );
  AOI22X1 U8486 ( .A0(n1187), .A1(x_matrix[26]), .B0(n1188), .B1(x_matrix[106]), .Y(n1275) );
  AOI22X1 U8487 ( .A0(n5298), .A1(x_matrix[186]), .B0(n5314), .B1(
        x_matrix[282]), .Y(n1274) );
  AOI221X1 U8488 ( .A0(n5289), .A1(x_matrix[554]), .B0(n5282), .B1(
        x_matrix[666]), .C0(n1277), .Y(n1276) );
  AOI31X1 U8489 ( .A0(n1539), .A1(n1540), .A2(n1541), .B0(n5318), .Y(N11594)
         );
  AOI22X1 U8490 ( .A0(n1455), .A1(x_matrix[618]), .B0(n1522), .B1(
        x_matrix[730]), .Y(n1539) );
  AOI22X1 U8491 ( .A0(n5258), .A1(x_matrix[410]), .B0(n5254), .B1(
        x_matrix[506]), .Y(n1540) );
  AOI221X1 U8492 ( .A0(n5295), .A1(x_matrix[218]), .B0(n5282), .B1(
        x_matrix[314]), .C0(n1542), .Y(n1541) );
  AOI31X1 U8493 ( .A0(n1270), .A1(n1271), .A2(n1272), .B0(n5321), .Y(N11975)
         );
  AOI22X1 U8494 ( .A0(n1187), .A1(x_matrix[27]), .B0(n1188), .B1(x_matrix[107]), .Y(n1271) );
  AOI22X1 U8495 ( .A0(n5298), .A1(x_matrix[187]), .B0(n5314), .B1(
        x_matrix[283]), .Y(n1270) );
  AOI221X1 U8496 ( .A0(n5291), .A1(x_matrix[555]), .B0(n5282), .B1(
        x_matrix[667]), .C0(n1273), .Y(n1272) );
  AOI31X1 U8497 ( .A0(n1535), .A1(n1536), .A2(n1537), .B0(n5318), .Y(N11595)
         );
  AOI22X1 U8498 ( .A0(n1455), .A1(x_matrix[619]), .B0(n1522), .B1(
        x_matrix[731]), .Y(n1535) );
  AOI22X1 U8499 ( .A0(n5257), .A1(x_matrix[411]), .B0(n5254), .B1(
        x_matrix[507]), .Y(n1536) );
  AOI221X1 U8500 ( .A0(n5295), .A1(x_matrix[219]), .B0(n5282), .B1(
        x_matrix[315]), .C0(n1538), .Y(n1537) );
  AOI31X1 U8501 ( .A0(n1266), .A1(n1267), .A2(n1268), .B0(n5321), .Y(N11976)
         );
  AOI22X1 U8502 ( .A0(n1187), .A1(x_matrix[28]), .B0(n1188), .B1(x_matrix[108]), .Y(n1267) );
  AOI22X1 U8503 ( .A0(n5298), .A1(x_matrix[188]), .B0(n5314), .B1(
        x_matrix[284]), .Y(n1266) );
  AOI221X1 U8504 ( .A0(n5291), .A1(x_matrix[556]), .B0(n5282), .B1(
        x_matrix[668]), .C0(n1269), .Y(n1268) );
  AOI31X1 U8505 ( .A0(n1531), .A1(n1532), .A2(n1533), .B0(n5318), .Y(N11596)
         );
  AOI22X1 U8506 ( .A0(n1455), .A1(x_matrix[620]), .B0(n1522), .B1(
        x_matrix[732]), .Y(n1531) );
  AOI22X1 U8507 ( .A0(n5257), .A1(x_matrix[412]), .B0(n5254), .B1(
        x_matrix[508]), .Y(n1532) );
  AOI221X1 U8508 ( .A0(n5294), .A1(x_matrix[220]), .B0(n5282), .B1(
        x_matrix[316]), .C0(n1534), .Y(n1533) );
  AOI31X1 U8509 ( .A0(n1262), .A1(n1263), .A2(n1264), .B0(n5321), .Y(N11977)
         );
  AOI22X1 U8510 ( .A0(n1187), .A1(x_matrix[29]), .B0(n1188), .B1(x_matrix[109]), .Y(n1263) );
  AOI22X1 U8511 ( .A0(n5298), .A1(x_matrix[189]), .B0(n5314), .B1(
        x_matrix[285]), .Y(n1262) );
  AOI221X1 U8512 ( .A0(n5289), .A1(x_matrix[557]), .B0(n5282), .B1(
        x_matrix[669]), .C0(n1265), .Y(n1264) );
  AOI31X1 U8513 ( .A0(n1527), .A1(n1528), .A2(n1529), .B0(n5318), .Y(N11597)
         );
  AOI22X1 U8514 ( .A0(n5251), .A1(x_matrix[621]), .B0(n1522), .B1(
        x_matrix[733]), .Y(n1527) );
  AOI22X1 U8515 ( .A0(n5257), .A1(x_matrix[413]), .B0(n1389), .B1(
        x_matrix[509]), .Y(n1528) );
  AOI221X1 U8516 ( .A0(n5294), .A1(x_matrix[221]), .B0(n5282), .B1(
        x_matrix[317]), .C0(n1530), .Y(n1529) );
  AOI31X1 U8517 ( .A0(n1238), .A1(n1239), .A2(n1240), .B0(n5321), .Y(N12062)
         );
  AOI22X1 U8518 ( .A0(n5060), .A1(x_matrix[2]), .B0(n1187), .B1(x_matrix[82]), 
        .Y(n1239) );
  AOI22X1 U8519 ( .A0(n5302), .A1(x_matrix[162]), .B0(n5299), .B1(
        x_matrix[258]), .Y(n1238) );
  AOI221X1 U8520 ( .A0(n5314), .A1(x_matrix[354]), .B0(n5272), .B1(
        x_matrix[450]), .C0(n1241), .Y(n1240) );
  AOI31X1 U8521 ( .A0(n1504), .A1(n1505), .A2(n1506), .B0(n5318), .Y(N11683)
         );
  AOI22X1 U8522 ( .A0(n5253), .A1(x_matrix[594]), .B0(n1455), .B1(
        x_matrix[706]), .Y(n1504) );
  AOI22X1 U8523 ( .A0(n5282), .A1(x_matrix[386]), .B0(n5258), .B1(
        x_matrix[482]), .Y(n1505) );
  AOI221X1 U8524 ( .A0(n1183), .A1(x_matrix[66]), .B0(n5277), .B1(
        x_matrix[146]), .C0(n1507), .Y(n1506) );
  AOI31X1 U8525 ( .A0(n1258), .A1(n1259), .A2(n1260), .B0(n5321), .Y(N11978)
         );
  AOI22X1 U8526 ( .A0(n1187), .A1(x_matrix[30]), .B0(n1188), .B1(x_matrix[110]), .Y(n1259) );
  AOI22X1 U8527 ( .A0(n5298), .A1(x_matrix[190]), .B0(n5314), .B1(
        x_matrix[286]), .Y(n1258) );
  AOI221X1 U8528 ( .A0(n5291), .A1(x_matrix[558]), .B0(n5282), .B1(
        x_matrix[670]), .C0(n1261), .Y(n1260) );
  AOI31X1 U8529 ( .A0(n1523), .A1(n1524), .A2(n1525), .B0(n5318), .Y(N11598)
         );
  AOI22X1 U8530 ( .A0(n1455), .A1(x_matrix[622]), .B0(n1522), .B1(
        x_matrix[734]), .Y(n1523) );
  AOI22X1 U8531 ( .A0(n5258), .A1(x_matrix[414]), .B0(n1389), .B1(
        x_matrix[510]), .Y(n1524) );
  AOI221X1 U8532 ( .A0(n5294), .A1(x_matrix[222]), .B0(n5282), .B1(
        x_matrix[318]), .C0(n1526), .Y(n1525) );
  AOI31X1 U8533 ( .A0(n1251), .A1(n1252), .A2(n1253), .B0(n5321), .Y(N11979)
         );
  AOI22X1 U8534 ( .A0(n1187), .A1(x_matrix[31]), .B0(n1188), .B1(x_matrix[111]), .Y(n1252) );
  AOI22X1 U8535 ( .A0(n5298), .A1(x_matrix[191]), .B0(n5314), .B1(
        x_matrix[287]), .Y(n1251) );
  AOI221X1 U8536 ( .A0(n5293), .A1(x_matrix[559]), .B0(n5282), .B1(
        x_matrix[671]), .C0(n1256), .Y(n1253) );
  AOI31X1 U8537 ( .A0(n1518), .A1(n1519), .A2(n1520), .B0(n5318), .Y(N11599)
         );
  AOI22X1 U8538 ( .A0(n1455), .A1(x_matrix[623]), .B0(n1522), .B1(
        x_matrix[735]), .Y(n1518) );
  AOI22X1 U8539 ( .A0(n5258), .A1(x_matrix[415]), .B0(n1389), .B1(
        x_matrix[511]), .Y(n1519) );
  AOI221X1 U8540 ( .A0(n5293), .A1(x_matrix[223]), .B0(n5282), .B1(
        x_matrix[319]), .C0(n1521), .Y(n1520) );
  AOI31X1 U8541 ( .A0(n1380), .A1(n1381), .A2(n1382), .B0(n5320), .Y(N11870)
         );
  AOI22X1 U8542 ( .A0(n5302), .A1(x_matrix[32]), .B0(n5299), .B1(x_matrix[112]), .Y(n1381) );
  AOI22X1 U8543 ( .A0(n1183), .A1(x_matrix[192]), .B0(n5265), .B1(
        x_matrix[288]), .Y(n1380) );
  AOI221X1 U8544 ( .A0(n5282), .A1(x_matrix[560]), .B0(n5257), .B1(
        x_matrix[672]), .C0(n1383), .Y(n1382) );
  AOI31X1 U8545 ( .A0(n1376), .A1(n1377), .A2(n1378), .B0(n5319), .Y(N11871)
         );
  AOI22X1 U8546 ( .A0(n5302), .A1(x_matrix[33]), .B0(n5299), .B1(x_matrix[113]), .Y(n1377) );
  AOI22X1 U8547 ( .A0(n1183), .A1(x_matrix[193]), .B0(n5267), .B1(
        x_matrix[289]), .Y(n1376) );
  AOI221X1 U8548 ( .A0(n5282), .A1(x_matrix[561]), .B0(n5257), .B1(
        x_matrix[673]), .C0(n1379), .Y(n1378) );
  AOI31X1 U8549 ( .A0(n1372), .A1(n1373), .A2(n1374), .B0(n5319), .Y(N11872)
         );
  AOI22X1 U8550 ( .A0(n1188), .A1(x_matrix[34]), .B0(n5299), .B1(x_matrix[114]), .Y(n1373) );
  AOI22X1 U8551 ( .A0(n1183), .A1(x_matrix[194]), .B0(n5270), .B1(
        x_matrix[290]), .Y(n1372) );
  AOI221X1 U8552 ( .A0(n5282), .A1(x_matrix[562]), .B0(n5257), .B1(
        x_matrix[674]), .C0(n1375), .Y(n1374) );
  AOI31X1 U8553 ( .A0(n1368), .A1(n1369), .A2(n1370), .B0(n5319), .Y(N11873)
         );
  AOI22X1 U8554 ( .A0(n5302), .A1(x_matrix[35]), .B0(n5299), .B1(x_matrix[115]), .Y(n1369) );
  AOI22X1 U8555 ( .A0(n1183), .A1(x_matrix[195]), .B0(n5266), .B1(
        x_matrix[291]), .Y(n1368) );
  AOI221X1 U8556 ( .A0(n5282), .A1(x_matrix[563]), .B0(n5257), .B1(
        x_matrix[675]), .C0(n1371), .Y(n1370) );
  AOI31X1 U8557 ( .A0(n1364), .A1(n1365), .A2(n1366), .B0(n5319), .Y(N11874)
         );
  AOI22X1 U8558 ( .A0(n1188), .A1(x_matrix[36]), .B0(n5299), .B1(x_matrix[116]), .Y(n1365) );
  AOI22X1 U8559 ( .A0(n1183), .A1(x_matrix[196]), .B0(n5272), .B1(
        x_matrix[292]), .Y(n1364) );
  AOI221X1 U8560 ( .A0(n5282), .A1(x_matrix[564]), .B0(n5259), .B1(
        x_matrix[676]), .C0(n1367), .Y(n1366) );
  AOI31X1 U8561 ( .A0(n1360), .A1(n1361), .A2(n1362), .B0(n5319), .Y(N11875)
         );
  AOI22X1 U8562 ( .A0(n5302), .A1(x_matrix[37]), .B0(n5299), .B1(x_matrix[117]), .Y(n1361) );
  AOI22X1 U8563 ( .A0(n1183), .A1(x_matrix[197]), .B0(n5267), .B1(
        x_matrix[293]), .Y(n1360) );
  AOI221X1 U8564 ( .A0(n5282), .A1(x_matrix[565]), .B0(n1322), .B1(
        x_matrix[677]), .C0(n1363), .Y(n1362) );
  AOI31X1 U8565 ( .A0(n1356), .A1(n1357), .A2(n1358), .B0(n5319), .Y(N11876)
         );
  AOI22X1 U8566 ( .A0(n1188), .A1(x_matrix[38]), .B0(n5299), .B1(x_matrix[118]), .Y(n1357) );
  AOI22X1 U8567 ( .A0(n1183), .A1(x_matrix[198]), .B0(n5265), .B1(
        x_matrix[294]), .Y(n1356) );
  AOI221X1 U8568 ( .A0(n5282), .A1(x_matrix[566]), .B0(n1322), .B1(
        x_matrix[678]), .C0(n1359), .Y(n1358) );
  AOI31X1 U8569 ( .A0(n1352), .A1(n1353), .A2(n1354), .B0(n5319), .Y(N11877)
         );
  AOI22X1 U8570 ( .A0(n5302), .A1(x_matrix[39]), .B0(n5299), .B1(x_matrix[119]), .Y(n1353) );
  AOI22X1 U8571 ( .A0(n1183), .A1(x_matrix[199]), .B0(n5268), .B1(
        x_matrix[295]), .Y(n1352) );
  AOI221X1 U8572 ( .A0(n5282), .A1(x_matrix[567]), .B0(n1322), .B1(
        x_matrix[679]), .C0(n1355), .Y(n1354) );
  AOI31X1 U8573 ( .A0(n1234), .A1(n1235), .A2(n1236), .B0(n5321), .Y(N12063)
         );
  AOI22X1 U8574 ( .A0(n5060), .A1(x_matrix[3]), .B0(n1187), .B1(x_matrix[83]), 
        .Y(n1235) );
  AOI22X1 U8575 ( .A0(n1188), .A1(x_matrix[163]), .B0(n1189), .B1(
        x_matrix[259]), .Y(n1234) );
  AOI221X1 U8576 ( .A0(n5314), .A1(x_matrix[355]), .B0(n5269), .B1(
        x_matrix[451]), .C0(n1237), .Y(n1236) );
  AOI31X1 U8577 ( .A0(n1500), .A1(n1501), .A2(n1502), .B0(n5318), .Y(N11684)
         );
  AOI22X1 U8578 ( .A0(n5253), .A1(x_matrix[595]), .B0(n1455), .B1(
        x_matrix[707]), .Y(n1500) );
  AOI22X1 U8579 ( .A0(n5282), .A1(x_matrix[387]), .B0(n5258), .B1(
        x_matrix[483]), .Y(n1501) );
  AOI221X1 U8580 ( .A0(n1183), .A1(x_matrix[67]), .B0(n5277), .B1(
        x_matrix[147]), .C0(n1503), .Y(n1502) );
  AOI31X1 U8581 ( .A0(n1348), .A1(n1349), .A2(n1350), .B0(n5319), .Y(N11878)
         );
  AOI22X1 U8582 ( .A0(n1188), .A1(x_matrix[40]), .B0(n5299), .B1(x_matrix[120]), .Y(n1349) );
  AOI22X1 U8583 ( .A0(n1183), .A1(x_matrix[200]), .B0(n5271), .B1(
        x_matrix[296]), .Y(n1348) );
  AOI221X1 U8584 ( .A0(n5282), .A1(x_matrix[568]), .B0(n1322), .B1(
        x_matrix[680]), .C0(n1351), .Y(n1350) );
  AOI31X1 U8585 ( .A0(n1344), .A1(n1345), .A2(n1346), .B0(n5319), .Y(N11879)
         );
  AOI22X1 U8586 ( .A0(n5302), .A1(x_matrix[41]), .B0(n1189), .B1(x_matrix[121]), .Y(n1345) );
  AOI22X1 U8587 ( .A0(n1183), .A1(x_matrix[201]), .B0(n5265), .B1(
        x_matrix[297]), .Y(n1344) );
  AOI221X1 U8588 ( .A0(n5282), .A1(x_matrix[569]), .B0(n1322), .B1(
        x_matrix[681]), .C0(n1347), .Y(n1346) );
  AOI31X1 U8589 ( .A0(n1340), .A1(n1341), .A2(n1342), .B0(n5319), .Y(N11880)
         );
  AOI22X1 U8590 ( .A0(n1188), .A1(x_matrix[42]), .B0(n5298), .B1(x_matrix[122]), .Y(n1341) );
  AOI22X1 U8591 ( .A0(n5314), .A1(x_matrix[202]), .B0(n5270), .B1(
        x_matrix[298]), .Y(n1340) );
  AOI221X1 U8592 ( .A0(n5282), .A1(x_matrix[570]), .B0(n1322), .B1(
        x_matrix[682]), .C0(n1343), .Y(n1342) );
  AOI31X1 U8593 ( .A0(n1336), .A1(n1337), .A2(n1338), .B0(n5319), .Y(N11881)
         );
  AOI22X1 U8594 ( .A0(n5302), .A1(x_matrix[43]), .B0(n1189), .B1(x_matrix[123]), .Y(n1337) );
  AOI22X1 U8595 ( .A0(n1183), .A1(x_matrix[203]), .B0(n5269), .B1(
        x_matrix[299]), .Y(n1336) );
  AOI221X1 U8596 ( .A0(n5282), .A1(x_matrix[571]), .B0(n1322), .B1(
        x_matrix[683]), .C0(n1339), .Y(n1338) );
  AOI31X1 U8597 ( .A0(n1332), .A1(n1333), .A2(n1334), .B0(n5319), .Y(N11882)
         );
  AOI22X1 U8598 ( .A0(n1188), .A1(x_matrix[44]), .B0(n5298), .B1(x_matrix[124]), .Y(n1333) );
  AOI22X1 U8599 ( .A0(n5314), .A1(x_matrix[204]), .B0(n5271), .B1(
        x_matrix[300]), .Y(n1332) );
  AOI221X1 U8600 ( .A0(n5282), .A1(x_matrix[572]), .B0(n1322), .B1(
        x_matrix[684]), .C0(n1335), .Y(n1334) );
  AOI31X1 U8601 ( .A0(n1328), .A1(n1329), .A2(n1330), .B0(n5319), .Y(N11883)
         );
  AOI22X1 U8602 ( .A0(n5302), .A1(x_matrix[45]), .B0(n1189), .B1(x_matrix[125]), .Y(n1329) );
  AOI22X1 U8603 ( .A0(n1183), .A1(x_matrix[205]), .B0(n5268), .B1(
        x_matrix[301]), .Y(n1328) );
  AOI221X1 U8604 ( .A0(n5282), .A1(x_matrix[573]), .B0(n1322), .B1(
        x_matrix[685]), .C0(n1331), .Y(n1330) );
  AOI31X1 U8605 ( .A0(n1324), .A1(n1325), .A2(n1326), .B0(n5320), .Y(N11884)
         );
  AOI22X1 U8606 ( .A0(n5302), .A1(x_matrix[46]), .B0(n5298), .B1(x_matrix[126]), .Y(n1325) );
  AOI22X1 U8607 ( .A0(n5314), .A1(x_matrix[206]), .B0(n5272), .B1(
        x_matrix[302]), .Y(n1324) );
  AOI221X1 U8608 ( .A0(n5282), .A1(x_matrix[574]), .B0(n1322), .B1(
        x_matrix[686]), .C0(n1327), .Y(n1326) );
  AOI31X1 U8609 ( .A0(n1319), .A1(n1320), .A2(n1321), .B0(n5320), .Y(N11885)
         );
  AOI22X1 U8610 ( .A0(n5302), .A1(x_matrix[47]), .B0(n1189), .B1(x_matrix[127]), .Y(n1320) );
  AOI22X1 U8611 ( .A0(n1183), .A1(x_matrix[207]), .B0(n5269), .B1(
        x_matrix[303]), .Y(n1319) );
  AOI221X1 U8612 ( .A0(n5282), .A1(x_matrix[575]), .B0(n1322), .B1(
        x_matrix[687]), .C0(n1323), .Y(n1321) );
  AOI31X1 U8613 ( .A0(n1446), .A1(n1447), .A2(n1448), .B0(n5317), .Y(N11773)
         );
  AOI22X1 U8614 ( .A0(n5293), .A1(x_matrix[368]), .B0(n5282), .B1(
        x_matrix[464]), .Y(n1447) );
  AOI22X1 U8615 ( .A0(n5257), .A1(x_matrix[576]), .B0(n1389), .B1(
        x_matrix[688]), .Y(n1446) );
  AOI221X1 U8616 ( .A0(n5299), .A1(x_matrix[48]), .B0(n5314), .B1(
        x_matrix[128]), .C0(n1449), .Y(n1448) );
  AOI31X1 U8617 ( .A0(n1442), .A1(n1443), .A2(n1444), .B0(n5318), .Y(N11774)
         );
  AOI22X1 U8618 ( .A0(n5290), .A1(x_matrix[369]), .B0(n5282), .B1(
        x_matrix[465]), .Y(n1443) );
  AOI22X1 U8619 ( .A0(n5258), .A1(x_matrix[577]), .B0(n1389), .B1(
        x_matrix[689]), .Y(n1442) );
  AOI221X1 U8620 ( .A0(n5299), .A1(x_matrix[49]), .B0(n5314), .B1(
        x_matrix[129]), .C0(n1445), .Y(n1444) );
  AOI31X1 U8621 ( .A0(n1230), .A1(n1231), .A2(n1232), .B0(n5321), .Y(N12064)
         );
  AOI22X1 U8622 ( .A0(n5060), .A1(x_matrix[4]), .B0(n1187), .B1(x_matrix[84]), 
        .Y(n1231) );
  AOI22X1 U8623 ( .A0(n1188), .A1(x_matrix[164]), .B0(n1189), .B1(
        x_matrix[260]), .Y(n1230) );
  AOI221X1 U8624 ( .A0(n5314), .A1(x_matrix[356]), .B0(n5272), .B1(
        x_matrix[452]), .C0(n1233), .Y(n1232) );
  AOI31X1 U8625 ( .A0(n1496), .A1(n1497), .A2(n1498), .B0(n5318), .Y(N11685)
         );
  AOI22X1 U8626 ( .A0(n5253), .A1(x_matrix[596]), .B0(n1455), .B1(
        x_matrix[708]), .Y(n1496) );
  AOI22X1 U8627 ( .A0(n5282), .A1(x_matrix[388]), .B0(n1322), .B1(
        x_matrix[484]), .Y(n1497) );
  AOI221X1 U8628 ( .A0(n1183), .A1(x_matrix[68]), .B0(n5277), .B1(
        x_matrix[148]), .C0(n1499), .Y(n1498) );
  AOI31X1 U8629 ( .A0(n1438), .A1(n1439), .A2(n1440), .B0(n5317), .Y(N11775)
         );
  AOI22X1 U8630 ( .A0(n5291), .A1(x_matrix[370]), .B0(n5282), .B1(
        x_matrix[466]), .Y(n1439) );
  AOI22X1 U8631 ( .A0(n1322), .A1(x_matrix[578]), .B0(n1389), .B1(
        x_matrix[690]), .Y(n1438) );
  AOI221X1 U8632 ( .A0(n5299), .A1(x_matrix[50]), .B0(n5314), .B1(
        x_matrix[130]), .C0(n1441), .Y(n1440) );
  AOI31X1 U8633 ( .A0(n1434), .A1(n1435), .A2(n1436), .B0(n5318), .Y(N11776)
         );
  AOI22X1 U8634 ( .A0(n5293), .A1(x_matrix[371]), .B0(n5282), .B1(
        x_matrix[467]), .Y(n1435) );
  AOI22X1 U8635 ( .A0(n5257), .A1(x_matrix[579]), .B0(n1389), .B1(
        x_matrix[691]), .Y(n1434) );
  AOI221X1 U8636 ( .A0(n5299), .A1(x_matrix[51]), .B0(n5314), .B1(
        x_matrix[131]), .C0(n1437), .Y(n1436) );
  AOI31X1 U8637 ( .A0(n1430), .A1(n1431), .A2(n1432), .B0(n5319), .Y(N11777)
         );
  AOI22X1 U8638 ( .A0(n5292), .A1(x_matrix[372]), .B0(n5282), .B1(
        x_matrix[468]), .Y(n1431) );
  AOI22X1 U8639 ( .A0(n1322), .A1(x_matrix[580]), .B0(n1389), .B1(
        x_matrix[692]), .Y(n1430) );
  AOI221X1 U8640 ( .A0(n5299), .A1(x_matrix[52]), .B0(n5314), .B1(
        x_matrix[132]), .C0(n1433), .Y(n1432) );
  AOI31X1 U8641 ( .A0(n1426), .A1(n1427), .A2(n1428), .B0(n5320), .Y(N11778)
         );
  AOI22X1 U8642 ( .A0(n5293), .A1(x_matrix[373]), .B0(n5282), .B1(
        x_matrix[469]), .Y(n1427) );
  AOI22X1 U8643 ( .A0(n5258), .A1(x_matrix[581]), .B0(n1389), .B1(
        x_matrix[693]), .Y(n1426) );
  AOI221X1 U8644 ( .A0(n5299), .A1(x_matrix[53]), .B0(n5314), .B1(
        x_matrix[133]), .C0(n1429), .Y(n1428) );
  AOI31X1 U8645 ( .A0(n1422), .A1(n1423), .A2(n1424), .B0(n5319), .Y(N11779)
         );
  AOI22X1 U8646 ( .A0(n5288), .A1(x_matrix[374]), .B0(n5282), .B1(
        x_matrix[470]), .Y(n1423) );
  AOI22X1 U8647 ( .A0(n1322), .A1(x_matrix[582]), .B0(n5254), .B1(
        x_matrix[694]), .Y(n1422) );
  AOI221X1 U8648 ( .A0(n5299), .A1(x_matrix[54]), .B0(n5314), .B1(
        x_matrix[134]), .C0(n1425), .Y(n1424) );
  AOI31X1 U8649 ( .A0(n1418), .A1(n1419), .A2(n1420), .B0(n5320), .Y(N11780)
         );
  AOI22X1 U8650 ( .A0(n5294), .A1(x_matrix[375]), .B0(n5282), .B1(
        x_matrix[471]), .Y(n1419) );
  AOI22X1 U8651 ( .A0(n5258), .A1(x_matrix[583]), .B0(n1389), .B1(
        x_matrix[695]), .Y(n1418) );
  AOI221X1 U8652 ( .A0(n5299), .A1(x_matrix[55]), .B0(n5314), .B1(
        x_matrix[135]), .C0(n1421), .Y(n1420) );
  AOI31X1 U8653 ( .A0(n1414), .A1(n1415), .A2(n1416), .B0(n5319), .Y(N11781)
         );
  AOI22X1 U8654 ( .A0(n5289), .A1(x_matrix[376]), .B0(n5282), .B1(
        x_matrix[472]), .Y(n1415) );
  AOI22X1 U8655 ( .A0(n1322), .A1(x_matrix[584]), .B0(n1389), .B1(
        x_matrix[696]), .Y(n1414) );
  AOI221X1 U8656 ( .A0(n5299), .A1(x_matrix[56]), .B0(n5314), .B1(
        x_matrix[136]), .C0(n1417), .Y(n1416) );
  AOI31X1 U8657 ( .A0(n1410), .A1(n1411), .A2(n1412), .B0(n5320), .Y(N11782)
         );
  AOI22X1 U8658 ( .A0(n5290), .A1(x_matrix[377]), .B0(n5282), .B1(
        x_matrix[473]), .Y(n1411) );
  AOI22X1 U8659 ( .A0(n5258), .A1(x_matrix[585]), .B0(n1389), .B1(
        x_matrix[697]), .Y(n1410) );
  AOI221X1 U8660 ( .A0(n5299), .A1(x_matrix[57]), .B0(n5314), .B1(
        x_matrix[137]), .C0(n1413), .Y(n1412) );
  AOI31X1 U8661 ( .A0(n1406), .A1(n1407), .A2(n1408), .B0(n5321), .Y(N11783)
         );
  AOI22X1 U8662 ( .A0(n5295), .A1(x_matrix[378]), .B0(n5282), .B1(
        x_matrix[474]), .Y(n1407) );
  AOI22X1 U8663 ( .A0(n5258), .A1(x_matrix[586]), .B0(n1389), .B1(
        x_matrix[698]), .Y(n1406) );
  AOI221X1 U8664 ( .A0(n5299), .A1(x_matrix[58]), .B0(n5314), .B1(
        x_matrix[138]), .C0(n1409), .Y(n1408) );
  AOI31X1 U8665 ( .A0(n1402), .A1(n1403), .A2(n1404), .B0(n5316), .Y(N11784)
         );
  AOI22X1 U8666 ( .A0(n5296), .A1(x_matrix[379]), .B0(n5282), .B1(
        x_matrix[475]), .Y(n1403) );
  AOI22X1 U8667 ( .A0(n5258), .A1(x_matrix[587]), .B0(n1389), .B1(
        x_matrix[699]), .Y(n1402) );
  AOI221X1 U8668 ( .A0(n5299), .A1(x_matrix[59]), .B0(n5314), .B1(
        x_matrix[139]), .C0(n1405), .Y(n1404) );
  AOI31X1 U8669 ( .A0(n1226), .A1(n1227), .A2(n1228), .B0(n5321), .Y(N12065)
         );
  AOI22X1 U8670 ( .A0(n5060), .A1(x_matrix[5]), .B0(n1187), .B1(x_matrix[85]), 
        .Y(n1227) );
  AOI22X1 U8671 ( .A0(n1188), .A1(x_matrix[165]), .B0(n1189), .B1(
        x_matrix[261]), .Y(n1226) );
  AOI221X1 U8672 ( .A0(n5314), .A1(x_matrix[357]), .B0(n5268), .B1(
        x_matrix[453]), .C0(n1229), .Y(n1228) );
  AOI31X1 U8673 ( .A0(n1492), .A1(n1493), .A2(n1494), .B0(n5318), .Y(N11686)
         );
  AOI22X1 U8674 ( .A0(n5253), .A1(x_matrix[597]), .B0(n1455), .B1(
        x_matrix[709]), .Y(n1492) );
  AOI22X1 U8675 ( .A0(n5282), .A1(x_matrix[389]), .B0(n1322), .B1(
        x_matrix[485]), .Y(n1493) );
  AOI221X1 U8676 ( .A0(n1183), .A1(x_matrix[69]), .B0(n5276), .B1(
        x_matrix[149]), .C0(n1495), .Y(n1494) );
  AOI31X1 U8677 ( .A0(n1398), .A1(n1399), .A2(n1400), .B0(n1182), .Y(N11785)
         );
  AOI22X1 U8678 ( .A0(n5292), .A1(x_matrix[380]), .B0(n5282), .B1(
        x_matrix[476]), .Y(n1399) );
  AOI22X1 U8679 ( .A0(n1322), .A1(x_matrix[588]), .B0(n1389), .B1(
        x_matrix[700]), .Y(n1398) );
  AOI221X1 U8680 ( .A0(n5299), .A1(x_matrix[60]), .B0(n5314), .B1(
        x_matrix[140]), .C0(n1401), .Y(n1400) );
  AOI31X1 U8681 ( .A0(n1394), .A1(n1395), .A2(n1396), .B0(n1182), .Y(N11786)
         );
  AOI22X1 U8682 ( .A0(n1254), .A1(x_matrix[381]), .B0(n5282), .B1(
        x_matrix[477]), .Y(n1395) );
  AOI22X1 U8683 ( .A0(n5258), .A1(x_matrix[589]), .B0(n1389), .B1(
        x_matrix[701]), .Y(n1394) );
  AOI221X1 U8684 ( .A0(n5299), .A1(x_matrix[61]), .B0(n5314), .B1(
        x_matrix[141]), .C0(n1397), .Y(n1396) );
  AOI31X1 U8685 ( .A0(n1390), .A1(n1391), .A2(n1392), .B0(n1182), .Y(N11787)
         );
  AOI22X1 U8686 ( .A0(n1254), .A1(x_matrix[382]), .B0(n5282), .B1(
        x_matrix[478]), .Y(n1391) );
  AOI22X1 U8687 ( .A0(n1322), .A1(x_matrix[590]), .B0(n1389), .B1(
        x_matrix[702]), .Y(n1390) );
  AOI221X1 U8688 ( .A0(n5299), .A1(x_matrix[62]), .B0(n5314), .B1(
        x_matrix[142]), .C0(n1393), .Y(n1392) );
  AOI31X1 U8689 ( .A0(n1385), .A1(n1386), .A2(n1387), .B0(n1182), .Y(N11788)
         );
  AOI22X1 U8690 ( .A0(n5294), .A1(x_matrix[383]), .B0(n5282), .B1(
        x_matrix[479]), .Y(n1386) );
  AOI22X1 U8691 ( .A0(n5257), .A1(x_matrix[591]), .B0(n1389), .B1(
        x_matrix[703]), .Y(n1385) );
  AOI221X1 U8692 ( .A0(n5299), .A1(x_matrix[63]), .B0(n5314), .B1(
        x_matrix[143]), .C0(n1388), .Y(n1387) );
  AOI31X1 U8693 ( .A0(n1222), .A1(n1223), .A2(n1224), .B0(n5321), .Y(N12066)
         );
  AOI22X1 U8694 ( .A0(n5060), .A1(x_matrix[6]), .B0(n1187), .B1(x_matrix[86]), 
        .Y(n1223) );
  AOI22X1 U8695 ( .A0(n1188), .A1(x_matrix[166]), .B0(n1189), .B1(
        x_matrix[262]), .Y(n1222) );
  AOI221X1 U8696 ( .A0(n5314), .A1(x_matrix[358]), .B0(n5270), .B1(
        x_matrix[454]), .C0(n1225), .Y(n1224) );
  AOI31X1 U8697 ( .A0(n1488), .A1(n1489), .A2(n1490), .B0(n5318), .Y(N11687)
         );
  AOI22X1 U8698 ( .A0(n5253), .A1(x_matrix[598]), .B0(n1455), .B1(
        x_matrix[710]), .Y(n1488) );
  AOI22X1 U8699 ( .A0(n5282), .A1(x_matrix[390]), .B0(n1322), .B1(
        x_matrix[486]), .Y(n1489) );
  AOI221X1 U8700 ( .A0(n1183), .A1(x_matrix[70]), .B0(n5276), .B1(
        x_matrix[150]), .C0(n1491), .Y(n1490) );
  AOI31X1 U8701 ( .A0(n1218), .A1(n1219), .A2(n1220), .B0(n5321), .Y(N12067)
         );
  AOI22X1 U8702 ( .A0(n5060), .A1(x_matrix[7]), .B0(n1187), .B1(x_matrix[87]), 
        .Y(n1219) );
  AOI22X1 U8703 ( .A0(n1188), .A1(x_matrix[167]), .B0(n1189), .B1(
        x_matrix[263]), .Y(n1218) );
  AOI221X1 U8704 ( .A0(n5314), .A1(x_matrix[359]), .B0(n5268), .B1(
        x_matrix[455]), .C0(n1221), .Y(n1220) );
  AOI31X1 U8705 ( .A0(n1484), .A1(n1485), .A2(n1486), .B0(n5319), .Y(N11688)
         );
  AOI22X1 U8706 ( .A0(n5253), .A1(x_matrix[599]), .B0(n1455), .B1(
        x_matrix[711]), .Y(n1484) );
  AOI22X1 U8707 ( .A0(n5282), .A1(x_matrix[391]), .B0(n1322), .B1(
        x_matrix[487]), .Y(n1485) );
  AOI221X1 U8708 ( .A0(n1183), .A1(x_matrix[71]), .B0(n5276), .B1(
        x_matrix[151]), .C0(n1487), .Y(n1486) );
  AOI31X1 U8709 ( .A0(n1480), .A1(n1481), .A2(n1482), .B0(n5320), .Y(N11689)
         );
  AOI22X1 U8710 ( .A0(n1389), .A1(x_matrix[600]), .B0(n1455), .B1(
        x_matrix[712]), .Y(n1480) );
  AOI22X1 U8711 ( .A0(n5282), .A1(x_matrix[392]), .B0(n1322), .B1(
        x_matrix[488]), .Y(n1481) );
  AOI221X1 U8712 ( .A0(n1183), .A1(x_matrix[72]), .B0(n5276), .B1(
        x_matrix[152]), .C0(n1483), .Y(n1482) );
  AOI31X1 U8713 ( .A0(n1476), .A1(n1477), .A2(n1478), .B0(n5319), .Y(N11690)
         );
  AOI22X1 U8714 ( .A0(n1389), .A1(x_matrix[601]), .B0(n1455), .B1(
        x_matrix[713]), .Y(n1476) );
  AOI22X1 U8715 ( .A0(n5282), .A1(x_matrix[393]), .B0(n1322), .B1(
        x_matrix[489]), .Y(n1477) );
  AOI221X1 U8716 ( .A0(n1183), .A1(x_matrix[73]), .B0(n5276), .B1(
        x_matrix[153]), .C0(n1479), .Y(n1478) );
  AND2X2 U8717 ( .A(N11313), .B(n1649), .Y(N11321) );
  AND2X2 U8718 ( .A(N11306), .B(n1649), .Y(N11314) );
  NOR3X1 U8719 ( .A(in_cnt_64[3]), .B(in_cnt_64[5]), .C(in_cnt_64[4]), .Y(
        n1517) );
  CLKINVX3 U8720 ( .A(c_plus[5]), .Y(n5935) );
  AND3X2 U8721 ( .A(in_addr_cnt[1]), .B(n4496), .C(n4497), .Y(n991) );
  OR3XL U8722 ( .A(mem_num_0), .B(n5064), .C(n5061), .Y(n4497) );
  CLKINVX3 U8723 ( .A(n1017), .Y(n5864) );
  AOI22X1 U8724 ( .A0(n5051), .A1(in_addr_cnt[4]), .B0(calweight_addr[4]), 
        .B1(n5066), .Y(n1017) );
  CLKINVX3 U8725 ( .A(n1025), .Y(n5872) );
  AOI22X1 U8726 ( .A0(n5051), .A1(in_addr_cnt[4]), .B0(calin_addr[4]), .B1(
        n5066), .Y(n1025) );
  CLKINVX3 U8727 ( .A(n1015), .Y(n5862) );
  AOI22X1 U8728 ( .A0(n5051), .A1(in_addr_cnt[6]), .B0(calweight_addr[6]), 
        .B1(n5066), .Y(n1015) );
  CLKINVX3 U8729 ( .A(n1023), .Y(n5870) );
  AOI22X1 U8730 ( .A0(n5051), .A1(in_addr_cnt[6]), .B0(calin_addr[6]), .B1(
        n5066), .Y(n1023) );
  CLKINVX3 U8731 ( .A(n1021), .Y(n5868) );
  AOI22X1 U8732 ( .A0(n5051), .A1(in_addr_cnt[0]), .B0(calweight_addr[0]), 
        .B1(n5066), .Y(n1021) );
  CLKINVX3 U8733 ( .A(n1029), .Y(n5876) );
  AOI22X1 U8734 ( .A0(n5051), .A1(in_addr_cnt[0]), .B0(calin_addr[0]), .B1(
        n5066), .Y(n1029) );
  OAI21XL U8735 ( .A0(N943), .A1(n746), .B0(n743), .Y(n742) );
  OAI22X1 U8736 ( .A0(n577), .A1(n5057), .B0(n625), .B1(n5058), .Y(n1717) );
  OAI22X1 U8737 ( .A0(n576), .A1(n5057), .B0(n624), .B1(n5058), .Y(n1713) );
  OAI22X1 U8738 ( .A0(n575), .A1(n5057), .B0(n623), .B1(n5058), .Y(n1709) );
  OAI22X1 U8739 ( .A0(n574), .A1(n5057), .B0(n622), .B1(n5058), .Y(n1705) );
  OAI22X1 U8740 ( .A0(n573), .A1(n5057), .B0(n621), .B1(n5058), .Y(n1701) );
  OAI22X1 U8741 ( .A0(n572), .A1(n5057), .B0(n620), .B1(n5058), .Y(n1697) );
  OAI22X1 U8742 ( .A0(n571), .A1(n5057), .B0(n619), .B1(n5058), .Y(n1693) );
  OAI22X1 U8743 ( .A0(n570), .A1(n5057), .B0(n618), .B1(n5058), .Y(n1689) );
  OAI22X1 U8744 ( .A0(n569), .A1(n5057), .B0(n617), .B1(n5058), .Y(n1685) );
  OAI22X1 U8745 ( .A0(n568), .A1(n5057), .B0(n616), .B1(n5058), .Y(n1681) );
  OAI22X1 U8746 ( .A0(n567), .A1(n5057), .B0(n615), .B1(n5058), .Y(n1677) );
  OAI22X1 U8747 ( .A0(n566), .A1(n5057), .B0(n614), .B1(n5058), .Y(n1673) );
  OAI22X1 U8748 ( .A0(n565), .A1(n5057), .B0(n613), .B1(n5058), .Y(n1669) );
  OAI22X1 U8749 ( .A0(n564), .A1(n5057), .B0(n612), .B1(n5058), .Y(n1665) );
  OAI22X1 U8750 ( .A0(n563), .A1(n5057), .B0(n611), .B1(n5058), .Y(n1661) );
  OAI22X1 U8751 ( .A0(n562), .A1(n5057), .B0(n610), .B1(n5058), .Y(n1657) );
  NAND3X1 U8752 ( .A(n828), .B(n5964), .C(c_plus[32]), .Y(n777) );
  NAND3X1 U8753 ( .A(n739), .B(n5051), .C(in_weight_flag), .Y(wen_weight) );
  NAND4X1 U8754 ( .A(n819), .B(n5931), .C(c_plus[0]), .D(n841), .Y(n840) );
  NOR3X1 U8755 ( .A(c_plus[35]), .B(c_plus[3]), .C(c_plus[37]), .Y(n841) );
  OR2X2 U8756 ( .A(out_cnt[1]), .B(out_cnt[0]), .Y(n5644) );
  AND3X2 U8757 ( .A(n803), .B(n5970), .C(n842), .Y(n819) );
  NOR3X1 U8758 ( .A(c_plus[4]), .B(c_plus[7]), .C(c_plus[5]), .Y(n842) );
  NAND3BX1 U8759 ( .AN(in_weight_flag), .B(n5052), .C(n739), .Y(wen_in) );
  OAI2BB2X1 U8760 ( .B0(n5939), .B1(n5596), .A0N(cal_out[9]), .A1N(n5189), .Y(
        n2402) );
  OAI2BB2X1 U8761 ( .B0(n5939), .B1(n5599), .A0N(cal_out[49]), .A1N(n5193), 
        .Y(n2362) );
  OAI2BB2X1 U8762 ( .B0(n5939), .B1(n5602), .A0N(cal_out[89]), .A1N(n5197), 
        .Y(n2322) );
  OAI2BB2X1 U8763 ( .B0(n5939), .B1(n5605), .A0N(cal_out[129]), .A1N(n5201), 
        .Y(n2282) );
  OAI2BB2X1 U8764 ( .B0(n5939), .B1(n5608), .A0N(cal_out[169]), .A1N(n5205), 
        .Y(n2242) );
  OAI2BB2X1 U8765 ( .B0(n5939), .B1(n5611), .A0N(cal_out[209]), .A1N(n5209), 
        .Y(n2202) );
  OAI2BB2X1 U8766 ( .B0(n5939), .B1(n5614), .A0N(cal_out[249]), .A1N(n5213), 
        .Y(n2162) );
  OAI2BB2X1 U8767 ( .B0(n5939), .B1(n5617), .A0N(cal_out[289]), .A1N(n5217), 
        .Y(n2122) );
  OAI2BB2X1 U8768 ( .B0(n5939), .B1(n5620), .A0N(cal_out[329]), .A1N(n5221), 
        .Y(n2082) );
  OAI2BB2X1 U8769 ( .B0(n5939), .B1(n5623), .A0N(cal_out[369]), .A1N(n5225), 
        .Y(n2042) );
  OAI2BB2X1 U8770 ( .B0(n5939), .B1(n5626), .A0N(cal_out[409]), .A1N(n5229), 
        .Y(n2002) );
  OAI2BB2XL U8771 ( .B0(n5939), .B1(n5629), .A0N(cal_out[449]), .A1N(n5233), 
        .Y(n1962) );
  OAI2BB2XL U8772 ( .B0(n5939), .B1(n5632), .A0N(cal_out[489]), .A1N(n5237), 
        .Y(n1922) );
  OAI2BB2XL U8773 ( .B0(n5939), .B1(n5634), .A0N(cal_out[529]), .A1N(n5856), 
        .Y(n1882) );
  OAI2BB2X1 U8774 ( .B0(n5950), .B1(n5596), .A0N(cal_out[19]), .A1N(n5190), 
        .Y(n2392) );
  OAI2BB2X1 U8775 ( .B0(n5950), .B1(n5599), .A0N(cal_out[59]), .A1N(n5194), 
        .Y(n2352) );
  OAI2BB2X1 U8776 ( .B0(n5950), .B1(n5602), .A0N(cal_out[99]), .A1N(n5198), 
        .Y(n2312) );
  OAI2BB2X1 U8777 ( .B0(n5950), .B1(n5605), .A0N(cal_out[139]), .A1N(n5202), 
        .Y(n2272) );
  OAI2BB2X1 U8778 ( .B0(n5950), .B1(n5608), .A0N(cal_out[179]), .A1N(n5206), 
        .Y(n2232) );
  OAI2BB2X1 U8779 ( .B0(n5950), .B1(n5611), .A0N(cal_out[219]), .A1N(n5210), 
        .Y(n2192) );
  OAI2BB2X1 U8780 ( .B0(n5950), .B1(n5614), .A0N(cal_out[259]), .A1N(n5214), 
        .Y(n2152) );
  OAI2BB2X1 U8781 ( .B0(n5950), .B1(n5617), .A0N(cal_out[299]), .A1N(n5218), 
        .Y(n2112) );
  OAI2BB2X1 U8782 ( .B0(n5950), .B1(n5620), .A0N(cal_out[339]), .A1N(n5222), 
        .Y(n2072) );
  OAI2BB2X1 U8783 ( .B0(n5950), .B1(n5623), .A0N(cal_out[379]), .A1N(n5226), 
        .Y(n2032) );
  OAI2BB2X1 U8784 ( .B0(n5950), .B1(n5626), .A0N(cal_out[419]), .A1N(n5230), 
        .Y(n1992) );
  OAI2BB2X1 U8785 ( .B0(n5950), .B1(n5629), .A0N(cal_out[459]), .A1N(n5234), 
        .Y(n1952) );
  OAI2BB2XL U8786 ( .B0(n5950), .B1(n5632), .A0N(cal_out[499]), .A1N(n5238), 
        .Y(n1912) );
  OAI2BB2XL U8787 ( .B0(n5950), .B1(n5634), .A0N(cal_out[539]), .A1N(n5241), 
        .Y(n1872) );
  OAI2BB2X1 U8788 ( .B0(n5954), .B1(n5595), .A0N(cal_out[23]), .A1N(n5190), 
        .Y(n2388) );
  OAI2BB2X1 U8789 ( .B0(n5954), .B1(n5598), .A0N(cal_out[63]), .A1N(n5194), 
        .Y(n2348) );
  OAI2BB2X1 U8790 ( .B0(n5954), .B1(n5601), .A0N(cal_out[103]), .A1N(n5198), 
        .Y(n2308) );
  OAI2BB2X1 U8791 ( .B0(n5954), .B1(n5604), .A0N(cal_out[143]), .A1N(n5202), 
        .Y(n2268) );
  OAI2BB2X1 U8792 ( .B0(n5954), .B1(n5607), .A0N(cal_out[183]), .A1N(n5206), 
        .Y(n2228) );
  OAI2BB2X1 U8793 ( .B0(n5954), .B1(n5610), .A0N(cal_out[223]), .A1N(n5210), 
        .Y(n2188) );
  OAI2BB2X1 U8794 ( .B0(n5954), .B1(n5613), .A0N(cal_out[263]), .A1N(n5214), 
        .Y(n2148) );
  OAI2BB2X1 U8795 ( .B0(n5954), .B1(n5616), .A0N(cal_out[303]), .A1N(n5218), 
        .Y(n2108) );
  OAI2BB2X1 U8796 ( .B0(n5954), .B1(n5619), .A0N(cal_out[343]), .A1N(n5222), 
        .Y(n2068) );
  OAI2BB2X1 U8797 ( .B0(n5954), .B1(n5622), .A0N(cal_out[383]), .A1N(n5226), 
        .Y(n2028) );
  OAI2BB2X1 U8798 ( .B0(n5954), .B1(n5625), .A0N(cal_out[423]), .A1N(n5230), 
        .Y(n1988) );
  OAI2BB2X1 U8799 ( .B0(n5954), .B1(n5628), .A0N(cal_out[463]), .A1N(n5234), 
        .Y(n1948) );
  OAI2BB2X1 U8800 ( .B0(n5954), .B1(n5631), .A0N(cal_out[503]), .A1N(n5238), 
        .Y(n1908) );
  OAI2BB2XL U8801 ( .B0(n5954), .B1(n5634), .A0N(cal_out[543]), .A1N(n5241), 
        .Y(n1868) );
  OAI2BB2X1 U8802 ( .B0(n5951), .B1(n5596), .A0N(cal_out[20]), .A1N(n5190), 
        .Y(n2391) );
  OAI2BB2X1 U8803 ( .B0(n5951), .B1(n5599), .A0N(cal_out[60]), .A1N(n5194), 
        .Y(n2351) );
  OAI2BB2X1 U8804 ( .B0(n5951), .B1(n5602), .A0N(cal_out[100]), .A1N(n5198), 
        .Y(n2311) );
  OAI2BB2X1 U8805 ( .B0(n5951), .B1(n5605), .A0N(cal_out[140]), .A1N(n5202), 
        .Y(n2271) );
  OAI2BB2X1 U8806 ( .B0(n5951), .B1(n5608), .A0N(cal_out[180]), .A1N(n5206), 
        .Y(n2231) );
  OAI2BB2X1 U8807 ( .B0(n5951), .B1(n5611), .A0N(cal_out[220]), .A1N(n5210), 
        .Y(n2191) );
  OAI2BB2X1 U8808 ( .B0(n5951), .B1(n5614), .A0N(cal_out[260]), .A1N(n5214), 
        .Y(n2151) );
  OAI2BB2X1 U8809 ( .B0(n5951), .B1(n5617), .A0N(cal_out[300]), .A1N(n5218), 
        .Y(n2111) );
  OAI2BB2X1 U8810 ( .B0(n5951), .B1(n5620), .A0N(cal_out[340]), .A1N(n5222), 
        .Y(n2071) );
  OAI2BB2X1 U8811 ( .B0(n5951), .B1(n5623), .A0N(cal_out[380]), .A1N(n5226), 
        .Y(n2031) );
  OAI2BB2X1 U8812 ( .B0(n5951), .B1(n5626), .A0N(cal_out[420]), .A1N(n5230), 
        .Y(n1991) );
  OAI2BB2X1 U8813 ( .B0(n5951), .B1(n5629), .A0N(cal_out[460]), .A1N(n5234), 
        .Y(n1951) );
  OAI2BB2X1 U8814 ( .B0(n5951), .B1(n5632), .A0N(cal_out[500]), .A1N(n5238), 
        .Y(n1911) );
  OAI2BB2XL U8815 ( .B0(n5951), .B1(n5634), .A0N(cal_out[540]), .A1N(n5241), 
        .Y(n1871) );
  OAI2BB2X1 U8816 ( .B0(n5959), .B1(n5595), .A0N(cal_out[27]), .A1N(n5191), 
        .Y(n2384) );
  OAI2BB2X1 U8817 ( .B0(n5959), .B1(n5598), .A0N(cal_out[67]), .A1N(n5195), 
        .Y(n2344) );
  OAI2BB2X1 U8818 ( .B0(n5959), .B1(n5601), .A0N(cal_out[107]), .A1N(n5199), 
        .Y(n2304) );
  OAI2BB2X1 U8819 ( .B0(n5959), .B1(n5604), .A0N(cal_out[147]), .A1N(n5203), 
        .Y(n2264) );
  OAI2BB2X1 U8820 ( .B0(n5959), .B1(n5607), .A0N(cal_out[187]), .A1N(n5207), 
        .Y(n2224) );
  OAI2BB2X1 U8821 ( .B0(n5959), .B1(n5610), .A0N(cal_out[227]), .A1N(n5211), 
        .Y(n2184) );
  OAI2BB2X1 U8822 ( .B0(n5959), .B1(n5613), .A0N(cal_out[267]), .A1N(n5215), 
        .Y(n2144) );
  OAI2BB2X1 U8823 ( .B0(n5959), .B1(n5616), .A0N(cal_out[307]), .A1N(n5219), 
        .Y(n2104) );
  OAI2BB2X1 U8824 ( .B0(n5959), .B1(n5619), .A0N(cal_out[347]), .A1N(n5223), 
        .Y(n2064) );
  OAI2BB2X1 U8825 ( .B0(n5959), .B1(n5622), .A0N(cal_out[387]), .A1N(n5227), 
        .Y(n2024) );
  OAI2BB2X1 U8826 ( .B0(n5959), .B1(n5625), .A0N(cal_out[427]), .A1N(n5231), 
        .Y(n1984) );
  OAI2BB2X1 U8827 ( .B0(n5959), .B1(n5628), .A0N(cal_out[467]), .A1N(n5235), 
        .Y(n1944) );
  OAI2BB2X1 U8828 ( .B0(n5959), .B1(n5631), .A0N(cal_out[507]), .A1N(n5239), 
        .Y(n1904) );
  OAI2BB2XL U8829 ( .B0(n5959), .B1(n5634), .A0N(cal_out[547]), .A1N(n5242), 
        .Y(n1864) );
  OAI2BB2X1 U8830 ( .B0(n5960), .B1(n5595), .A0N(cal_out[28]), .A1N(n5191), 
        .Y(n2383) );
  OAI2BB2X1 U8831 ( .B0(n5960), .B1(n5598), .A0N(cal_out[68]), .A1N(n5195), 
        .Y(n2343) );
  OAI2BB2X1 U8832 ( .B0(n5960), .B1(n5601), .A0N(cal_out[108]), .A1N(n5199), 
        .Y(n2303) );
  OAI2BB2X1 U8833 ( .B0(n5960), .B1(n5604), .A0N(cal_out[148]), .A1N(n5203), 
        .Y(n2263) );
  OAI2BB2X1 U8834 ( .B0(n5960), .B1(n5607), .A0N(cal_out[188]), .A1N(n5207), 
        .Y(n2223) );
  OAI2BB2X1 U8835 ( .B0(n5960), .B1(n5610), .A0N(cal_out[228]), .A1N(n5211), 
        .Y(n2183) );
  OAI2BB2X1 U8836 ( .B0(n5960), .B1(n5613), .A0N(cal_out[268]), .A1N(n5215), 
        .Y(n2143) );
  OAI2BB2X1 U8837 ( .B0(n5960), .B1(n5616), .A0N(cal_out[308]), .A1N(n5219), 
        .Y(n2103) );
  OAI2BB2X1 U8838 ( .B0(n5960), .B1(n5619), .A0N(cal_out[348]), .A1N(n5223), 
        .Y(n2063) );
  OAI2BB2X1 U8839 ( .B0(n5960), .B1(n5622), .A0N(cal_out[388]), .A1N(n5227), 
        .Y(n2023) );
  OAI2BB2X1 U8840 ( .B0(n5960), .B1(n5625), .A0N(cal_out[428]), .A1N(n5231), 
        .Y(n1983) );
  OAI2BB2X1 U8841 ( .B0(n5960), .B1(n5628), .A0N(cal_out[468]), .A1N(n5235), 
        .Y(n1943) );
  OAI2BB2X1 U8842 ( .B0(n5960), .B1(n5631), .A0N(cal_out[508]), .A1N(n5239), 
        .Y(n1903) );
  OAI2BB2XL U8843 ( .B0(n5960), .B1(n5634), .A0N(cal_out[548]), .A1N(n5242), 
        .Y(n1863) );
  OAI2BB2X1 U8844 ( .B0(n5953), .B1(n5595), .A0N(cal_out[22]), .A1N(n5190), 
        .Y(n2389) );
  OAI2BB2X1 U8845 ( .B0(n5953), .B1(n5598), .A0N(cal_out[62]), .A1N(n5194), 
        .Y(n2349) );
  OAI2BB2X1 U8846 ( .B0(n5953), .B1(n5601), .A0N(cal_out[102]), .A1N(n5198), 
        .Y(n2309) );
  OAI2BB2X1 U8847 ( .B0(n5953), .B1(n5604), .A0N(cal_out[142]), .A1N(n5202), 
        .Y(n2269) );
  OAI2BB2X1 U8848 ( .B0(n5953), .B1(n5607), .A0N(cal_out[182]), .A1N(n5206), 
        .Y(n2229) );
  OAI2BB2X1 U8849 ( .B0(n5953), .B1(n5610), .A0N(cal_out[222]), .A1N(n5210), 
        .Y(n2189) );
  OAI2BB2X1 U8850 ( .B0(n5953), .B1(n5613), .A0N(cal_out[262]), .A1N(n5214), 
        .Y(n2149) );
  OAI2BB2X1 U8851 ( .B0(n5953), .B1(n5616), .A0N(cal_out[302]), .A1N(n5218), 
        .Y(n2109) );
  OAI2BB2X1 U8852 ( .B0(n5953), .B1(n5619), .A0N(cal_out[342]), .A1N(n5222), 
        .Y(n2069) );
  OAI2BB2X1 U8853 ( .B0(n5953), .B1(n5622), .A0N(cal_out[382]), .A1N(n5226), 
        .Y(n2029) );
  OAI2BB2X1 U8854 ( .B0(n5953), .B1(n5625), .A0N(cal_out[422]), .A1N(n5230), 
        .Y(n1989) );
  OAI2BB2X1 U8855 ( .B0(n5953), .B1(n5628), .A0N(cal_out[462]), .A1N(n5234), 
        .Y(n1949) );
  OAI2BB2X1 U8856 ( .B0(n5953), .B1(n5631), .A0N(cal_out[502]), .A1N(n5238), 
        .Y(n1909) );
  OAI2BB2XL U8857 ( .B0(n5953), .B1(n5634), .A0N(cal_out[542]), .A1N(n5241), 
        .Y(n1869) );
  OAI2BB2X1 U8858 ( .B0(n5935), .B1(n5596), .A0N(cal_out[5]), .A1N(n5189), .Y(
        n2406) );
  OAI2BB2X1 U8859 ( .B0(n5935), .B1(n5599), .A0N(cal_out[45]), .A1N(n5193), 
        .Y(n2366) );
  OAI2BB2X1 U8860 ( .B0(n5935), .B1(n5602), .A0N(cal_out[85]), .A1N(n5197), 
        .Y(n2326) );
  OAI2BB2X1 U8861 ( .B0(n5935), .B1(n5605), .A0N(cal_out[125]), .A1N(n5201), 
        .Y(n2286) );
  OAI2BB2X1 U8862 ( .B0(n5935), .B1(n5608), .A0N(cal_out[165]), .A1N(n5205), 
        .Y(n2246) );
  OAI2BB2X1 U8863 ( .B0(n5935), .B1(n5611), .A0N(cal_out[205]), .A1N(n5209), 
        .Y(n2206) );
  OAI2BB2X1 U8864 ( .B0(n5935), .B1(n5614), .A0N(cal_out[245]), .A1N(n5213), 
        .Y(n2166) );
  OAI2BB2X1 U8865 ( .B0(n5935), .B1(n5617), .A0N(cal_out[285]), .A1N(n5217), 
        .Y(n2126) );
  OAI2BB2X1 U8866 ( .B0(n5935), .B1(n5620), .A0N(cal_out[325]), .A1N(n5221), 
        .Y(n2086) );
  OAI2BB2X1 U8867 ( .B0(n5935), .B1(n5623), .A0N(cal_out[365]), .A1N(n5225), 
        .Y(n2046) );
  OAI2BB2X1 U8868 ( .B0(n5935), .B1(n5626), .A0N(cal_out[405]), .A1N(n5229), 
        .Y(n2006) );
  OAI2BB2X1 U8869 ( .B0(n5935), .B1(n5629), .A0N(cal_out[445]), .A1N(n5233), 
        .Y(n1966) );
  OAI2BB2X1 U8870 ( .B0(n5935), .B1(n5632), .A0N(cal_out[485]), .A1N(n5237), 
        .Y(n1926) );
  OAI2BB2XL U8871 ( .B0(n5935), .B1(n5635), .A0N(cal_out[525]), .A1N(n5856), 
        .Y(n1886) );
  OAI2BB2X1 U8872 ( .B0(n5965), .B1(n5594), .A0N(cal_out[34]), .A1N(n5191), 
        .Y(n2377) );
  OAI2BB2X1 U8873 ( .B0(n5965), .B1(n5597), .A0N(cal_out[74]), .A1N(n5195), 
        .Y(n2337) );
  OAI2BB2X1 U8874 ( .B0(n5965), .B1(n5600), .A0N(cal_out[114]), .A1N(n5199), 
        .Y(n2297) );
  OAI2BB2X1 U8875 ( .B0(n5965), .B1(n5603), .A0N(cal_out[154]), .A1N(n5203), 
        .Y(n2257) );
  OAI2BB2X1 U8876 ( .B0(n5965), .B1(n5606), .A0N(cal_out[194]), .A1N(n5207), 
        .Y(n2217) );
  OAI2BB2X1 U8877 ( .B0(n5965), .B1(n5609), .A0N(cal_out[234]), .A1N(n5211), 
        .Y(n2177) );
  OAI2BB2X1 U8878 ( .B0(n5965), .B1(n5612), .A0N(cal_out[274]), .A1N(n5215), 
        .Y(n2137) );
  OAI2BB2X1 U8879 ( .B0(n5965), .B1(n5615), .A0N(cal_out[314]), .A1N(n5219), 
        .Y(n2097) );
  OAI2BB2X1 U8880 ( .B0(n5965), .B1(n5618), .A0N(cal_out[354]), .A1N(n5223), 
        .Y(n2057) );
  OAI2BB2X1 U8881 ( .B0(n5965), .B1(n5621), .A0N(cal_out[394]), .A1N(n5227), 
        .Y(n2017) );
  OAI2BB2X1 U8882 ( .B0(n5965), .B1(n5624), .A0N(cal_out[434]), .A1N(n5231), 
        .Y(n1977) );
  OAI2BB2X1 U8883 ( .B0(n5965), .B1(n5627), .A0N(cal_out[474]), .A1N(n5235), 
        .Y(n1937) );
  OAI2BB2X1 U8884 ( .B0(n5965), .B1(n5630), .A0N(cal_out[514]), .A1N(n5239), 
        .Y(n1897) );
  OAI2BB2XL U8885 ( .B0(n5965), .B1(n5633), .A0N(cal_out[554]), .A1N(n5242), 
        .Y(n1857) );
  OAI2BB2XL U8886 ( .B0(n5965), .B1(n5637), .A0N(cal_out[594]), .A1N(n5247), 
        .Y(n1817) );
  OAI2BB2X1 U8887 ( .B0(n5934), .B1(n5596), .A0N(cal_out[4]), .A1N(n5189), .Y(
        n2407) );
  OAI2BB2X1 U8888 ( .B0(n5934), .B1(n5599), .A0N(cal_out[44]), .A1N(n5193), 
        .Y(n2367) );
  OAI2BB2X1 U8889 ( .B0(n5934), .B1(n5602), .A0N(cal_out[84]), .A1N(n5197), 
        .Y(n2327) );
  OAI2BB2X1 U8890 ( .B0(n5934), .B1(n5605), .A0N(cal_out[124]), .A1N(n5201), 
        .Y(n2287) );
  OAI2BB2X1 U8891 ( .B0(n5934), .B1(n5608), .A0N(cal_out[164]), .A1N(n5205), 
        .Y(n2247) );
  OAI2BB2X1 U8892 ( .B0(n5934), .B1(n5611), .A0N(cal_out[204]), .A1N(n5209), 
        .Y(n2207) );
  OAI2BB2X1 U8893 ( .B0(n5934), .B1(n5614), .A0N(cal_out[244]), .A1N(n5213), 
        .Y(n2167) );
  OAI2BB2X1 U8894 ( .B0(n5934), .B1(n5617), .A0N(cal_out[284]), .A1N(n5217), 
        .Y(n2127) );
  OAI2BB2X1 U8895 ( .B0(n5934), .B1(n5620), .A0N(cal_out[324]), .A1N(n5221), 
        .Y(n2087) );
  OAI2BB2X1 U8896 ( .B0(n5934), .B1(n5623), .A0N(cal_out[364]), .A1N(n5225), 
        .Y(n2047) );
  OAI2BB2X1 U8897 ( .B0(n5934), .B1(n5626), .A0N(cal_out[404]), .A1N(n5229), 
        .Y(n2007) );
  OAI2BB2X1 U8898 ( .B0(n5934), .B1(n5629), .A0N(cal_out[444]), .A1N(n5233), 
        .Y(n1967) );
  OAI2BB2X1 U8899 ( .B0(n5934), .B1(n5632), .A0N(cal_out[484]), .A1N(n5237), 
        .Y(n1927) );
  OAI2BB2X1 U8900 ( .B0(n5934), .B1(n5635), .A0N(cal_out[524]), .A1N(n5243), 
        .Y(n1887) );
  OAI2BB2X1 U8901 ( .B0(n5957), .B1(n5595), .A0N(cal_out[25]), .A1N(n5191), 
        .Y(n2386) );
  OAI2BB2X1 U8902 ( .B0(n5957), .B1(n5598), .A0N(cal_out[65]), .A1N(n5195), 
        .Y(n2346) );
  OAI2BB2X1 U8903 ( .B0(n5957), .B1(n5601), .A0N(cal_out[105]), .A1N(n5199), 
        .Y(n2306) );
  OAI2BB2X1 U8904 ( .B0(n5957), .B1(n5604), .A0N(cal_out[145]), .A1N(n5203), 
        .Y(n2266) );
  OAI2BB2X1 U8905 ( .B0(n5957), .B1(n5607), .A0N(cal_out[185]), .A1N(n5207), 
        .Y(n2226) );
  OAI2BB2X1 U8906 ( .B0(n5957), .B1(n5610), .A0N(cal_out[225]), .A1N(n5211), 
        .Y(n2186) );
  OAI2BB2X1 U8907 ( .B0(n5957), .B1(n5613), .A0N(cal_out[265]), .A1N(n5215), 
        .Y(n2146) );
  OAI2BB2X1 U8908 ( .B0(n5957), .B1(n5616), .A0N(cal_out[305]), .A1N(n5219), 
        .Y(n2106) );
  OAI2BB2X1 U8909 ( .B0(n5957), .B1(n5619), .A0N(cal_out[345]), .A1N(n5223), 
        .Y(n2066) );
  OAI2BB2X1 U8910 ( .B0(n5957), .B1(n5622), .A0N(cal_out[385]), .A1N(n5227), 
        .Y(n2026) );
  OAI2BB2X1 U8911 ( .B0(n5957), .B1(n5625), .A0N(cal_out[425]), .A1N(n5231), 
        .Y(n1986) );
  OAI2BB2X1 U8912 ( .B0(n5957), .B1(n5628), .A0N(cal_out[465]), .A1N(n5235), 
        .Y(n1946) );
  OAI2BB2XL U8913 ( .B0(n5957), .B1(n5631), .A0N(cal_out[505]), .A1N(n5239), 
        .Y(n1906) );
  OAI2BB2XL U8914 ( .B0(n5957), .B1(n5634), .A0N(cal_out[545]), .A1N(n5242), 
        .Y(n1866) );
  OAI2BB2X1 U8915 ( .B0(n5944), .B1(n5596), .A0N(cal_out[13]), .A1N(n5190), 
        .Y(n2398) );
  OAI2BB2X1 U8916 ( .B0(n5944), .B1(n5599), .A0N(cal_out[53]), .A1N(n5194), 
        .Y(n2358) );
  OAI2BB2X1 U8917 ( .B0(n5944), .B1(n5602), .A0N(cal_out[93]), .A1N(n5198), 
        .Y(n2318) );
  OAI2BB2X1 U8918 ( .B0(n5944), .B1(n5605), .A0N(cal_out[133]), .A1N(n5202), 
        .Y(n2278) );
  OAI2BB2X1 U8919 ( .B0(n5944), .B1(n5608), .A0N(cal_out[173]), .A1N(n5206), 
        .Y(n2238) );
  OAI2BB2X1 U8920 ( .B0(n5944), .B1(n5611), .A0N(cal_out[213]), .A1N(n5210), 
        .Y(n2198) );
  OAI2BB2X1 U8921 ( .B0(n5944), .B1(n5614), .A0N(cal_out[253]), .A1N(n5214), 
        .Y(n2158) );
  OAI2BB2X1 U8922 ( .B0(n5944), .B1(n5617), .A0N(cal_out[293]), .A1N(n5218), 
        .Y(n2118) );
  OAI2BB2X1 U8923 ( .B0(n5944), .B1(n5620), .A0N(cal_out[333]), .A1N(n5222), 
        .Y(n2078) );
  OAI2BB2X1 U8924 ( .B0(n5944), .B1(n5623), .A0N(cal_out[373]), .A1N(n5226), 
        .Y(n2038) );
  OAI2BB2X1 U8925 ( .B0(n5944), .B1(n5626), .A0N(cal_out[413]), .A1N(n5230), 
        .Y(n1998) );
  OAI2BB2X1 U8926 ( .B0(n5944), .B1(n5629), .A0N(cal_out[453]), .A1N(n5234), 
        .Y(n1958) );
  OAI2BB2X1 U8927 ( .B0(n5944), .B1(n5632), .A0N(cal_out[493]), .A1N(n5238), 
        .Y(n1918) );
  OAI2BB2XL U8928 ( .B0(n5944), .B1(n5634), .A0N(cal_out[533]), .A1N(n5241), 
        .Y(n1878) );
  OAI2BB2X1 U8929 ( .B0(n5938), .B1(n5596), .A0N(cal_out[8]), .A1N(n5189), .Y(
        n2403) );
  OAI2BB2X1 U8930 ( .B0(n5938), .B1(n5599), .A0N(cal_out[48]), .A1N(n5193), 
        .Y(n2363) );
  OAI2BB2X1 U8931 ( .B0(n5938), .B1(n5602), .A0N(cal_out[88]), .A1N(n5197), 
        .Y(n2323) );
  OAI2BB2X1 U8932 ( .B0(n5938), .B1(n5605), .A0N(cal_out[128]), .A1N(n5201), 
        .Y(n2283) );
  OAI2BB2X1 U8933 ( .B0(n5938), .B1(n5608), .A0N(cal_out[168]), .A1N(n5205), 
        .Y(n2243) );
  OAI2BB2X1 U8934 ( .B0(n5938), .B1(n5611), .A0N(cal_out[208]), .A1N(n5209), 
        .Y(n2203) );
  OAI2BB2X1 U8935 ( .B0(n5938), .B1(n5614), .A0N(cal_out[248]), .A1N(n5213), 
        .Y(n2163) );
  OAI2BB2X1 U8936 ( .B0(n5938), .B1(n5617), .A0N(cal_out[288]), .A1N(n5217), 
        .Y(n2123) );
  OAI2BB2X1 U8937 ( .B0(n5938), .B1(n5620), .A0N(cal_out[328]), .A1N(n5221), 
        .Y(n2083) );
  OAI2BB2X1 U8938 ( .B0(n5938), .B1(n5623), .A0N(cal_out[368]), .A1N(n5225), 
        .Y(n2043) );
  OAI2BB2X1 U8939 ( .B0(n5938), .B1(n5626), .A0N(cal_out[408]), .A1N(n5229), 
        .Y(n2003) );
  OAI2BB2X1 U8940 ( .B0(n5938), .B1(n5629), .A0N(cal_out[448]), .A1N(n5233), 
        .Y(n1963) );
  OAI2BB2XL U8941 ( .B0(n5938), .B1(n5632), .A0N(cal_out[488]), .A1N(n5237), 
        .Y(n1923) );
  OAI2BB2XL U8942 ( .B0(n5938), .B1(n5634), .A0N(cal_out[528]), .A1N(n5856), 
        .Y(n1883) );
  OAI2BB2X1 U8943 ( .B0(n5931), .B1(n5595), .A0N(cal_out[1]), .A1N(n5189), .Y(
        n2410) );
  OAI2BB2X1 U8944 ( .B0(n5931), .B1(n5598), .A0N(cal_out[41]), .A1N(n5193), 
        .Y(n2370) );
  OAI2BB2X1 U8945 ( .B0(n5931), .B1(n5601), .A0N(cal_out[81]), .A1N(n5197), 
        .Y(n2330) );
  OAI2BB2X1 U8946 ( .B0(n5931), .B1(n5604), .A0N(cal_out[121]), .A1N(n5201), 
        .Y(n2290) );
  OAI2BB2X1 U8947 ( .B0(n5931), .B1(n5607), .A0N(cal_out[161]), .A1N(n5205), 
        .Y(n2250) );
  OAI2BB2X1 U8948 ( .B0(n5931), .B1(n5610), .A0N(cal_out[201]), .A1N(n5209), 
        .Y(n2210) );
  OAI2BB2X1 U8949 ( .B0(n5931), .B1(n5613), .A0N(cal_out[241]), .A1N(n5213), 
        .Y(n2170) );
  OAI2BB2X1 U8950 ( .B0(n5931), .B1(n5616), .A0N(cal_out[281]), .A1N(n5217), 
        .Y(n2130) );
  OAI2BB2X1 U8951 ( .B0(n5931), .B1(n5619), .A0N(cal_out[321]), .A1N(n5221), 
        .Y(n2090) );
  OAI2BB2X1 U8952 ( .B0(n5931), .B1(n5622), .A0N(cal_out[361]), .A1N(n5225), 
        .Y(n2050) );
  OAI2BB2X1 U8953 ( .B0(n5931), .B1(n5625), .A0N(cal_out[401]), .A1N(n5229), 
        .Y(n2010) );
  OAI2BB2X1 U8954 ( .B0(n5931), .B1(n5628), .A0N(cal_out[441]), .A1N(n5233), 
        .Y(n1970) );
  OAI2BB2XL U8955 ( .B0(n5931), .B1(n5632), .A0N(cal_out[481]), .A1N(n5237), 
        .Y(n1930) );
  OAI2BB2XL U8956 ( .B0(n5931), .B1(n5635), .A0N(cal_out[521]), .A1N(n5856), 
        .Y(n1890) );
  OAI2BB2X1 U8957 ( .B0(n5961), .B1(n5595), .A0N(cal_out[29]), .A1N(n5191), 
        .Y(n2382) );
  OAI2BB2X1 U8958 ( .B0(n5961), .B1(n5598), .A0N(cal_out[69]), .A1N(n5195), 
        .Y(n2342) );
  OAI2BB2X1 U8959 ( .B0(n5961), .B1(n5601), .A0N(cal_out[109]), .A1N(n5199), 
        .Y(n2302) );
  OAI2BB2X1 U8960 ( .B0(n5961), .B1(n5604), .A0N(cal_out[149]), .A1N(n5203), 
        .Y(n2262) );
  OAI2BB2X1 U8961 ( .B0(n5961), .B1(n5607), .A0N(cal_out[189]), .A1N(n5207), 
        .Y(n2222) );
  OAI2BB2X1 U8962 ( .B0(n5961), .B1(n5610), .A0N(cal_out[229]), .A1N(n5211), 
        .Y(n2182) );
  OAI2BB2X1 U8963 ( .B0(n5961), .B1(n5613), .A0N(cal_out[269]), .A1N(n5215), 
        .Y(n2142) );
  OAI2BB2X1 U8964 ( .B0(n5961), .B1(n5616), .A0N(cal_out[309]), .A1N(n5219), 
        .Y(n2102) );
  OAI2BB2X1 U8965 ( .B0(n5961), .B1(n5619), .A0N(cal_out[349]), .A1N(n5223), 
        .Y(n2062) );
  OAI2BB2X1 U8966 ( .B0(n5961), .B1(n5622), .A0N(cal_out[389]), .A1N(n5227), 
        .Y(n2022) );
  OAI2BB2X1 U8967 ( .B0(n5961), .B1(n5625), .A0N(cal_out[429]), .A1N(n5231), 
        .Y(n1982) );
  OAI2BB2X1 U8968 ( .B0(n5961), .B1(n5628), .A0N(cal_out[469]), .A1N(n5235), 
        .Y(n1942) );
  OAI2BB2XL U8969 ( .B0(n5961), .B1(n5631), .A0N(cal_out[509]), .A1N(n5239), 
        .Y(n1902) );
  OAI2BB2XL U8970 ( .B0(n5961), .B1(n5633), .A0N(cal_out[549]), .A1N(n5242), 
        .Y(n1862) );
  OAI2BB2X1 U8971 ( .B0(n5958), .B1(n5595), .A0N(cal_out[26]), .A1N(n5191), 
        .Y(n2385) );
  OAI2BB2X1 U8972 ( .B0(n5958), .B1(n5598), .A0N(cal_out[66]), .A1N(n5195), 
        .Y(n2345) );
  OAI2BB2X1 U8973 ( .B0(n5958), .B1(n5601), .A0N(cal_out[106]), .A1N(n5199), 
        .Y(n2305) );
  OAI2BB2X1 U8974 ( .B0(n5958), .B1(n5604), .A0N(cal_out[146]), .A1N(n5203), 
        .Y(n2265) );
  OAI2BB2X1 U8975 ( .B0(n5958), .B1(n5607), .A0N(cal_out[186]), .A1N(n5207), 
        .Y(n2225) );
  OAI2BB2X1 U8976 ( .B0(n5958), .B1(n5610), .A0N(cal_out[226]), .A1N(n5211), 
        .Y(n2185) );
  OAI2BB2X1 U8977 ( .B0(n5958), .B1(n5613), .A0N(cal_out[266]), .A1N(n5215), 
        .Y(n2145) );
  OAI2BB2X1 U8978 ( .B0(n5958), .B1(n5616), .A0N(cal_out[306]), .A1N(n5219), 
        .Y(n2105) );
  OAI2BB2X1 U8979 ( .B0(n5958), .B1(n5619), .A0N(cal_out[346]), .A1N(n5223), 
        .Y(n2065) );
  OAI2BB2X1 U8980 ( .B0(n5958), .B1(n5622), .A0N(cal_out[386]), .A1N(n5227), 
        .Y(n2025) );
  OAI2BB2X1 U8981 ( .B0(n5958), .B1(n5625), .A0N(cal_out[426]), .A1N(n5231), 
        .Y(n1985) );
  OAI2BB2X1 U8982 ( .B0(n5958), .B1(n5628), .A0N(cal_out[466]), .A1N(n5235), 
        .Y(n1945) );
  OAI2BB2XL U8983 ( .B0(n5958), .B1(n5631), .A0N(cal_out[506]), .A1N(n5239), 
        .Y(n1905) );
  OAI2BB2XL U8984 ( .B0(n5958), .B1(n5633), .A0N(cal_out[546]), .A1N(n5242), 
        .Y(n1865) );
  OAI2BB2X1 U8985 ( .B0(n5955), .B1(n5595), .A0N(cal_out[24]), .A1N(n5191), 
        .Y(n2387) );
  OAI2BB2X1 U8986 ( .B0(n5955), .B1(n5598), .A0N(cal_out[64]), .A1N(n5195), 
        .Y(n2347) );
  OAI2BB2X1 U8987 ( .B0(n5955), .B1(n5601), .A0N(cal_out[104]), .A1N(n5199), 
        .Y(n2307) );
  OAI2BB2X1 U8988 ( .B0(n5955), .B1(n5604), .A0N(cal_out[144]), .A1N(n5203), 
        .Y(n2267) );
  OAI2BB2X1 U8989 ( .B0(n5955), .B1(n5607), .A0N(cal_out[184]), .A1N(n5207), 
        .Y(n2227) );
  OAI2BB2X1 U8990 ( .B0(n5955), .B1(n5610), .A0N(cal_out[224]), .A1N(n5211), 
        .Y(n2187) );
  OAI2BB2X1 U8991 ( .B0(n5955), .B1(n5613), .A0N(cal_out[264]), .A1N(n5215), 
        .Y(n2147) );
  OAI2BB2X1 U8992 ( .B0(n5955), .B1(n5616), .A0N(cal_out[304]), .A1N(n5219), 
        .Y(n2107) );
  OAI2BB2X1 U8993 ( .B0(n5955), .B1(n5619), .A0N(cal_out[344]), .A1N(n5223), 
        .Y(n2067) );
  OAI2BB2X1 U8994 ( .B0(n5955), .B1(n5622), .A0N(cal_out[384]), .A1N(n5227), 
        .Y(n2027) );
  OAI2BB2X1 U8995 ( .B0(n5955), .B1(n5625), .A0N(cal_out[424]), .A1N(n5231), 
        .Y(n1987) );
  OAI2BB2X1 U8996 ( .B0(n5955), .B1(n5628), .A0N(cal_out[464]), .A1N(n5235), 
        .Y(n1947) );
  OAI2BB2XL U8997 ( .B0(n5955), .B1(n5631), .A0N(cal_out[504]), .A1N(n5239), 
        .Y(n1907) );
  OAI2BB2XL U8998 ( .B0(n5955), .B1(n5634), .A0N(cal_out[544]), .A1N(n5242), 
        .Y(n1867) );
  OAI2BB2X1 U8999 ( .B0(n5967), .B1(n5594), .A0N(cal_out[36]), .A1N(n5843), 
        .Y(n2375) );
  OAI2BB2X1 U9000 ( .B0(n5967), .B1(n5597), .A0N(cal_out[76]), .A1N(n5844), 
        .Y(n2335) );
  OAI2BB2X1 U9001 ( .B0(n5967), .B1(n5600), .A0N(cal_out[116]), .A1N(n5845), 
        .Y(n2295) );
  OAI2BB2X1 U9002 ( .B0(n5967), .B1(n5603), .A0N(cal_out[156]), .A1N(n5846), 
        .Y(n2255) );
  OAI2BB2X1 U9003 ( .B0(n5967), .B1(n5606), .A0N(cal_out[196]), .A1N(n5847), 
        .Y(n2215) );
  OAI2BB2X1 U9004 ( .B0(n5967), .B1(n5609), .A0N(cal_out[236]), .A1N(n5848), 
        .Y(n2175) );
  OAI2BB2X1 U9005 ( .B0(n5967), .B1(n5612), .A0N(cal_out[276]), .A1N(n5849), 
        .Y(n2135) );
  OAI2BB2X1 U9006 ( .B0(n5967), .B1(n5615), .A0N(cal_out[316]), .A1N(n5850), 
        .Y(n2095) );
  OAI2BB2X1 U9007 ( .B0(n5967), .B1(n5618), .A0N(cal_out[356]), .A1N(n5851), 
        .Y(n2055) );
  OAI2BB2X1 U9008 ( .B0(n5967), .B1(n5621), .A0N(cal_out[396]), .A1N(n5852), 
        .Y(n2015) );
  OAI2BB2X1 U9009 ( .B0(n5967), .B1(n5624), .A0N(cal_out[436]), .A1N(n5853), 
        .Y(n1975) );
  OAI2BB2X1 U9010 ( .B0(n5967), .B1(n5627), .A0N(cal_out[476]), .A1N(n5854), 
        .Y(n1935) );
  OAI2BB2XL U9011 ( .B0(n5967), .B1(n5630), .A0N(cal_out[516]), .A1N(n5855), 
        .Y(n1895) );
  OAI2BB2XL U9012 ( .B0(n5967), .B1(n5633), .A0N(cal_out[556]), .A1N(n5243), 
        .Y(n1855) );
  OAI2BB2XL U9013 ( .B0(n5967), .B1(n5637), .A0N(cal_out[596]), .A1N(n5857), 
        .Y(n1815) );
  OAI2BB2X1 U9014 ( .B0(n5963), .B1(n5595), .A0N(cal_out[32]), .A1N(n5191), 
        .Y(n2379) );
  OAI2BB2X1 U9015 ( .B0(n5963), .B1(n5598), .A0N(cal_out[72]), .A1N(n5195), 
        .Y(n2339) );
  OAI2BB2X1 U9016 ( .B0(n5963), .B1(n5601), .A0N(cal_out[112]), .A1N(n5199), 
        .Y(n2299) );
  OAI2BB2X1 U9017 ( .B0(n5963), .B1(n5604), .A0N(cal_out[152]), .A1N(n5203), 
        .Y(n2259) );
  OAI2BB2X1 U9018 ( .B0(n5963), .B1(n5607), .A0N(cal_out[192]), .A1N(n5207), 
        .Y(n2219) );
  OAI2BB2X1 U9019 ( .B0(n5963), .B1(n5610), .A0N(cal_out[232]), .A1N(n5211), 
        .Y(n2179) );
  OAI2BB2X1 U9020 ( .B0(n5963), .B1(n5613), .A0N(cal_out[272]), .A1N(n5215), 
        .Y(n2139) );
  OAI2BB2X1 U9021 ( .B0(n5963), .B1(n5616), .A0N(cal_out[312]), .A1N(n5219), 
        .Y(n2099) );
  OAI2BB2X1 U9022 ( .B0(n5963), .B1(n5619), .A0N(cal_out[352]), .A1N(n5223), 
        .Y(n2059) );
  OAI2BB2X1 U9023 ( .B0(n5963), .B1(n5622), .A0N(cal_out[392]), .A1N(n5227), 
        .Y(n2019) );
  OAI2BB2X1 U9024 ( .B0(n5963), .B1(n5625), .A0N(cal_out[432]), .A1N(n5231), 
        .Y(n1979) );
  OAI2BB2X1 U9025 ( .B0(n5963), .B1(n5628), .A0N(cal_out[472]), .A1N(n5235), 
        .Y(n1939) );
  OAI2BB2XL U9026 ( .B0(n5963), .B1(n5631), .A0N(cal_out[512]), .A1N(n5239), 
        .Y(n1899) );
  OAI2BB2XL U9027 ( .B0(n5963), .B1(n5633), .A0N(cal_out[552]), .A1N(n5242), 
        .Y(n1859) );
  OAI2BB2XL U9028 ( .B0(n5963), .B1(n5637), .A0N(cal_out[592]), .A1N(n5247), 
        .Y(n1819) );
  OAI2BB2X1 U9029 ( .B0(n5946), .B1(n5596), .A0N(cal_out[15]), .A1N(n5190), 
        .Y(n2396) );
  OAI2BB2X1 U9030 ( .B0(n5946), .B1(n5599), .A0N(cal_out[55]), .A1N(n5194), 
        .Y(n2356) );
  OAI2BB2X1 U9031 ( .B0(n5946), .B1(n5602), .A0N(cal_out[95]), .A1N(n5198), 
        .Y(n2316) );
  OAI2BB2X1 U9032 ( .B0(n5946), .B1(n5605), .A0N(cal_out[135]), .A1N(n5202), 
        .Y(n2276) );
  OAI2BB2X1 U9033 ( .B0(n5946), .B1(n5608), .A0N(cal_out[175]), .A1N(n5206), 
        .Y(n2236) );
  OAI2BB2X1 U9034 ( .B0(n5946), .B1(n5611), .A0N(cal_out[215]), .A1N(n5210), 
        .Y(n2196) );
  OAI2BB2X1 U9035 ( .B0(n5946), .B1(n5614), .A0N(cal_out[255]), .A1N(n5214), 
        .Y(n2156) );
  OAI2BB2X1 U9036 ( .B0(n5946), .B1(n5617), .A0N(cal_out[295]), .A1N(n5218), 
        .Y(n2116) );
  OAI2BB2X1 U9037 ( .B0(n5946), .B1(n5620), .A0N(cal_out[335]), .A1N(n5222), 
        .Y(n2076) );
  OAI2BB2X1 U9038 ( .B0(n5946), .B1(n5623), .A0N(cal_out[375]), .A1N(n5226), 
        .Y(n2036) );
  OAI2BB2X1 U9039 ( .B0(n5946), .B1(n5626), .A0N(cal_out[415]), .A1N(n5230), 
        .Y(n1996) );
  OAI2BB2X1 U9040 ( .B0(n5946), .B1(n5629), .A0N(cal_out[455]), .A1N(n5234), 
        .Y(n1956) );
  OAI2BB2X1 U9041 ( .B0(n5946), .B1(n5632), .A0N(cal_out[495]), .A1N(n5238), 
        .Y(n1916) );
  OAI2BB2X1 U9042 ( .B0(n5946), .B1(n5634), .A0N(cal_out[535]), .A1N(n5241), 
        .Y(n1876) );
  OAI2BB2X1 U9043 ( .B0(n5942), .B1(n5596), .A0N(cal_out[11]), .A1N(n5189), 
        .Y(n2400) );
  OAI2BB2X1 U9044 ( .B0(n5942), .B1(n5599), .A0N(cal_out[51]), .A1N(n5193), 
        .Y(n2360) );
  OAI2BB2X1 U9045 ( .B0(n5942), .B1(n5602), .A0N(cal_out[91]), .A1N(n5197), 
        .Y(n2320) );
  OAI2BB2X1 U9046 ( .B0(n5942), .B1(n5605), .A0N(cal_out[131]), .A1N(n5201), 
        .Y(n2280) );
  OAI2BB2X1 U9047 ( .B0(n5942), .B1(n5608), .A0N(cal_out[171]), .A1N(n5205), 
        .Y(n2240) );
  OAI2BB2X1 U9048 ( .B0(n5942), .B1(n5611), .A0N(cal_out[211]), .A1N(n5209), 
        .Y(n2200) );
  OAI2BB2X1 U9049 ( .B0(n5942), .B1(n5614), .A0N(cal_out[251]), .A1N(n5213), 
        .Y(n2160) );
  OAI2BB2X1 U9050 ( .B0(n5942), .B1(n5617), .A0N(cal_out[291]), .A1N(n5217), 
        .Y(n2120) );
  OAI2BB2X1 U9051 ( .B0(n5942), .B1(n5620), .A0N(cal_out[331]), .A1N(n5221), 
        .Y(n2080) );
  OAI2BB2X1 U9052 ( .B0(n5942), .B1(n5623), .A0N(cal_out[371]), .A1N(n5225), 
        .Y(n2040) );
  OAI2BB2X1 U9053 ( .B0(n5942), .B1(n5626), .A0N(cal_out[411]), .A1N(n5229), 
        .Y(n2000) );
  OAI2BB2X1 U9054 ( .B0(n5942), .B1(n5629), .A0N(cal_out[451]), .A1N(n5233), 
        .Y(n1960) );
  OAI2BB2XL U9055 ( .B0(n5942), .B1(n5632), .A0N(cal_out[491]), .A1N(n5237), 
        .Y(n1920) );
  OAI2BB2XL U9056 ( .B0(n5942), .B1(n5634), .A0N(cal_out[531]), .A1N(n5856), 
        .Y(n1880) );
  OAI2BB2X1 U9057 ( .B0(n5947), .B1(n5596), .A0N(cal_out[16]), .A1N(n5190), 
        .Y(n2395) );
  OAI2BB2X1 U9058 ( .B0(n5947), .B1(n5599), .A0N(cal_out[56]), .A1N(n5194), 
        .Y(n2355) );
  OAI2BB2X1 U9059 ( .B0(n5947), .B1(n5602), .A0N(cal_out[96]), .A1N(n5198), 
        .Y(n2315) );
  OAI2BB2X1 U9060 ( .B0(n5947), .B1(n5605), .A0N(cal_out[136]), .A1N(n5202), 
        .Y(n2275) );
  OAI2BB2X1 U9061 ( .B0(n5947), .B1(n5608), .A0N(cal_out[176]), .A1N(n5206), 
        .Y(n2235) );
  OAI2BB2X1 U9062 ( .B0(n5947), .B1(n5611), .A0N(cal_out[216]), .A1N(n5210), 
        .Y(n2195) );
  OAI2BB2X1 U9063 ( .B0(n5947), .B1(n5614), .A0N(cal_out[256]), .A1N(n5214), 
        .Y(n2155) );
  OAI2BB2X1 U9064 ( .B0(n5947), .B1(n5617), .A0N(cal_out[296]), .A1N(n5218), 
        .Y(n2115) );
  OAI2BB2X1 U9065 ( .B0(n5947), .B1(n5620), .A0N(cal_out[336]), .A1N(n5222), 
        .Y(n2075) );
  OAI2BB2X1 U9066 ( .B0(n5947), .B1(n5623), .A0N(cal_out[376]), .A1N(n5226), 
        .Y(n2035) );
  OAI2BB2X1 U9067 ( .B0(n5947), .B1(n5626), .A0N(cal_out[416]), .A1N(n5230), 
        .Y(n1995) );
  OAI2BB2X1 U9068 ( .B0(n5947), .B1(n5629), .A0N(cal_out[456]), .A1N(n5234), 
        .Y(n1955) );
  OAI2BB2X1 U9069 ( .B0(n5947), .B1(n5632), .A0N(cal_out[496]), .A1N(n5238), 
        .Y(n1915) );
  OAI2BB2X1 U9070 ( .B0(n5947), .B1(n5634), .A0N(cal_out[536]), .A1N(n5241), 
        .Y(n1875) );
  OAI2BB2X1 U9071 ( .B0(n5940), .B1(n5596), .A0N(cal_out[10]), .A1N(n5189), 
        .Y(n2401) );
  OAI2BB2X1 U9072 ( .B0(n5940), .B1(n5599), .A0N(cal_out[50]), .A1N(n5193), 
        .Y(n2361) );
  OAI2BB2X1 U9073 ( .B0(n5940), .B1(n5602), .A0N(cal_out[90]), .A1N(n5197), 
        .Y(n2321) );
  OAI2BB2X1 U9074 ( .B0(n5940), .B1(n5605), .A0N(cal_out[130]), .A1N(n5201), 
        .Y(n2281) );
  OAI2BB2X1 U9075 ( .B0(n5940), .B1(n5608), .A0N(cal_out[170]), .A1N(n5205), 
        .Y(n2241) );
  OAI2BB2X1 U9076 ( .B0(n5940), .B1(n5611), .A0N(cal_out[210]), .A1N(n5209), 
        .Y(n2201) );
  OAI2BB2X1 U9077 ( .B0(n5940), .B1(n5614), .A0N(cal_out[250]), .A1N(n5213), 
        .Y(n2161) );
  OAI2BB2X1 U9078 ( .B0(n5940), .B1(n5617), .A0N(cal_out[290]), .A1N(n5217), 
        .Y(n2121) );
  OAI2BB2X1 U9079 ( .B0(n5940), .B1(n5620), .A0N(cal_out[330]), .A1N(n5221), 
        .Y(n2081) );
  OAI2BB2X1 U9080 ( .B0(n5940), .B1(n5623), .A0N(cal_out[370]), .A1N(n5225), 
        .Y(n2041) );
  OAI2BB2X1 U9081 ( .B0(n5940), .B1(n5626), .A0N(cal_out[410]), .A1N(n5229), 
        .Y(n2001) );
  OAI2BB2X1 U9082 ( .B0(n5940), .B1(n5629), .A0N(cal_out[450]), .A1N(n5233), 
        .Y(n1961) );
  OAI2BB2X1 U9083 ( .B0(n5940), .B1(n5632), .A0N(cal_out[490]), .A1N(n5237), 
        .Y(n1921) );
  OAI2BB2XL U9084 ( .B0(n5940), .B1(n5634), .A0N(cal_out[530]), .A1N(n5856), 
        .Y(n1881) );
  OAI2BB2X1 U9085 ( .B0(n5949), .B1(n5596), .A0N(cal_out[18]), .A1N(n5190), 
        .Y(n2393) );
  OAI2BB2X1 U9086 ( .B0(n5949), .B1(n5599), .A0N(cal_out[58]), .A1N(n5194), 
        .Y(n2353) );
  OAI2BB2X1 U9087 ( .B0(n5949), .B1(n5602), .A0N(cal_out[98]), .A1N(n5198), 
        .Y(n2313) );
  OAI2BB2X1 U9088 ( .B0(n5949), .B1(n5605), .A0N(cal_out[138]), .A1N(n5202), 
        .Y(n2273) );
  OAI2BB2X1 U9089 ( .B0(n5949), .B1(n5608), .A0N(cal_out[178]), .A1N(n5206), 
        .Y(n2233) );
  OAI2BB2X1 U9090 ( .B0(n5949), .B1(n5611), .A0N(cal_out[218]), .A1N(n5210), 
        .Y(n2193) );
  OAI2BB2X1 U9091 ( .B0(n5949), .B1(n5614), .A0N(cal_out[258]), .A1N(n5214), 
        .Y(n2153) );
  OAI2BB2X1 U9092 ( .B0(n5949), .B1(n5617), .A0N(cal_out[298]), .A1N(n5218), 
        .Y(n2113) );
  OAI2BB2X1 U9093 ( .B0(n5949), .B1(n5620), .A0N(cal_out[338]), .A1N(n5222), 
        .Y(n2073) );
  OAI2BB2X1 U9094 ( .B0(n5949), .B1(n5623), .A0N(cal_out[378]), .A1N(n5226), 
        .Y(n2033) );
  OAI2BB2X1 U9095 ( .B0(n5949), .B1(n5626), .A0N(cal_out[418]), .A1N(n5230), 
        .Y(n1993) );
  OAI2BB2X1 U9096 ( .B0(n5949), .B1(n5629), .A0N(cal_out[458]), .A1N(n5234), 
        .Y(n1953) );
  OAI2BB2X1 U9097 ( .B0(n5949), .B1(n5632), .A0N(cal_out[498]), .A1N(n5238), 
        .Y(n1913) );
  OAI2BB2XL U9098 ( .B0(n5949), .B1(n5634), .A0N(cal_out[538]), .A1N(n5241), 
        .Y(n1873) );
  OAI2BB2X1 U9099 ( .B0(n5937), .B1(n5596), .A0N(cal_out[7]), .A1N(n5189), .Y(
        n2404) );
  OAI2BB2X1 U9100 ( .B0(n5937), .B1(n5599), .A0N(cal_out[47]), .A1N(n5193), 
        .Y(n2364) );
  OAI2BB2X1 U9101 ( .B0(n5937), .B1(n5602), .A0N(cal_out[87]), .A1N(n5197), 
        .Y(n2324) );
  OAI2BB2X1 U9102 ( .B0(n5937), .B1(n5605), .A0N(cal_out[127]), .A1N(n5201), 
        .Y(n2284) );
  OAI2BB2X1 U9103 ( .B0(n5937), .B1(n5608), .A0N(cal_out[167]), .A1N(n5205), 
        .Y(n2244) );
  OAI2BB2X1 U9104 ( .B0(n5937), .B1(n5611), .A0N(cal_out[207]), .A1N(n5209), 
        .Y(n2204) );
  OAI2BB2X1 U9105 ( .B0(n5937), .B1(n5614), .A0N(cal_out[247]), .A1N(n5213), 
        .Y(n2164) );
  OAI2BB2X1 U9106 ( .B0(n5937), .B1(n5617), .A0N(cal_out[287]), .A1N(n5217), 
        .Y(n2124) );
  OAI2BB2X1 U9107 ( .B0(n5937), .B1(n5620), .A0N(cal_out[327]), .A1N(n5221), 
        .Y(n2084) );
  OAI2BB2X1 U9108 ( .B0(n5937), .B1(n5623), .A0N(cal_out[367]), .A1N(n5225), 
        .Y(n2044) );
  OAI2BB2X1 U9109 ( .B0(n5937), .B1(n5626), .A0N(cal_out[407]), .A1N(n5229), 
        .Y(n2004) );
  OAI2BB2X1 U9110 ( .B0(n5937), .B1(n5629), .A0N(cal_out[447]), .A1N(n5233), 
        .Y(n1964) );
  OAI2BB2X1 U9111 ( .B0(n5937), .B1(n5632), .A0N(cal_out[487]), .A1N(n5237), 
        .Y(n1924) );
  OAI2BB2XL U9112 ( .B0(n5937), .B1(n5635), .A0N(cal_out[527]), .A1N(n5856), 
        .Y(n1884) );
  NAND2X1 U9113 ( .A(c_plus[34]), .B(n854), .Y(n782) );
  OAI2BB2X1 U9114 ( .B0(n5943), .B1(n5596), .A0N(cal_out[12]), .A1N(n5190), 
        .Y(n2399) );
  OAI2BB2X1 U9115 ( .B0(n5943), .B1(n5599), .A0N(cal_out[52]), .A1N(n5194), 
        .Y(n2359) );
  OAI2BB2X1 U9116 ( .B0(n5943), .B1(n5602), .A0N(cal_out[92]), .A1N(n5198), 
        .Y(n2319) );
  OAI2BB2X1 U9117 ( .B0(n5943), .B1(n5605), .A0N(cal_out[132]), .A1N(n5202), 
        .Y(n2279) );
  OAI2BB2X1 U9118 ( .B0(n5943), .B1(n5608), .A0N(cal_out[172]), .A1N(n5206), 
        .Y(n2239) );
  OAI2BB2X1 U9119 ( .B0(n5943), .B1(n5611), .A0N(cal_out[212]), .A1N(n5210), 
        .Y(n2199) );
  OAI2BB2X1 U9120 ( .B0(n5943), .B1(n5614), .A0N(cal_out[252]), .A1N(n5214), 
        .Y(n2159) );
  OAI2BB2X1 U9121 ( .B0(n5943), .B1(n5617), .A0N(cal_out[292]), .A1N(n5218), 
        .Y(n2119) );
  OAI2BB2X1 U9122 ( .B0(n5943), .B1(n5620), .A0N(cal_out[332]), .A1N(n5222), 
        .Y(n2079) );
  OAI2BB2X1 U9123 ( .B0(n5943), .B1(n5623), .A0N(cal_out[372]), .A1N(n5226), 
        .Y(n2039) );
  OAI2BB2X1 U9124 ( .B0(n5943), .B1(n5626), .A0N(cal_out[412]), .A1N(n5230), 
        .Y(n1999) );
  OAI2BB2X1 U9125 ( .B0(n5943), .B1(n5629), .A0N(cal_out[452]), .A1N(n5234), 
        .Y(n1959) );
  OAI2BB2X1 U9126 ( .B0(n5943), .B1(n5632), .A0N(cal_out[492]), .A1N(n5238), 
        .Y(n1919) );
  OAI2BB2XL U9127 ( .B0(n5943), .B1(n5634), .A0N(cal_out[532]), .A1N(n5241), 
        .Y(n1879) );
  OAI2BB2X1 U9128 ( .B0(n5930), .B1(n5594), .A0N(cal_out[0]), .A1N(n5189), .Y(
        n2411) );
  OAI2BB2X1 U9129 ( .B0(n5930), .B1(n5597), .A0N(cal_out[40]), .A1N(n5193), 
        .Y(n2371) );
  OAI2BB2X1 U9130 ( .B0(n5930), .B1(n5600), .A0N(cal_out[80]), .A1N(n5197), 
        .Y(n2331) );
  OAI2BB2X1 U9131 ( .B0(n5930), .B1(n5603), .A0N(cal_out[120]), .A1N(n5201), 
        .Y(n2291) );
  OAI2BB2X1 U9132 ( .B0(n5930), .B1(n5606), .A0N(cal_out[160]), .A1N(n5205), 
        .Y(n2251) );
  OAI2BB2X1 U9133 ( .B0(n5930), .B1(n5609), .A0N(cal_out[200]), .A1N(n5209), 
        .Y(n2211) );
  OAI2BB2X1 U9134 ( .B0(n5930), .B1(n5612), .A0N(cal_out[240]), .A1N(n5213), 
        .Y(n2171) );
  OAI2BB2X1 U9135 ( .B0(n5930), .B1(n5615), .A0N(cal_out[280]), .A1N(n5217), 
        .Y(n2131) );
  OAI2BB2X1 U9136 ( .B0(n5930), .B1(n5618), .A0N(cal_out[320]), .A1N(n5221), 
        .Y(n2091) );
  OAI2BB2X1 U9137 ( .B0(n5930), .B1(n5621), .A0N(cal_out[360]), .A1N(n5225), 
        .Y(n2051) );
  OAI2BB2X1 U9138 ( .B0(n5930), .B1(n5624), .A0N(cal_out[400]), .A1N(n5229), 
        .Y(n2011) );
  OAI2BB2X1 U9139 ( .B0(n5930), .B1(n5627), .A0N(cal_out[440]), .A1N(n5233), 
        .Y(n1971) );
  OAI2BB2X1 U9140 ( .B0(n5930), .B1(n5630), .A0N(cal_out[480]), .A1N(n5237), 
        .Y(n1931) );
  OAI2BB2X1 U9141 ( .B0(n5930), .B1(n5633), .A0N(cal_out[520]), .A1N(n5856), 
        .Y(n1891) );
  OAI2BB2X1 U9142 ( .B0(n5936), .B1(n5594), .A0N(cal_out[6]), .A1N(n5189), .Y(
        n2405) );
  OAI2BB2X1 U9143 ( .B0(n5936), .B1(n5597), .A0N(cal_out[46]), .A1N(n5193), 
        .Y(n2365) );
  OAI2BB2X1 U9144 ( .B0(n5936), .B1(n5600), .A0N(cal_out[86]), .A1N(n5197), 
        .Y(n2325) );
  OAI2BB2X1 U9145 ( .B0(n5936), .B1(n5603), .A0N(cal_out[126]), .A1N(n5201), 
        .Y(n2285) );
  OAI2BB2X1 U9146 ( .B0(n5936), .B1(n5606), .A0N(cal_out[166]), .A1N(n5205), 
        .Y(n2245) );
  OAI2BB2X1 U9147 ( .B0(n5936), .B1(n5609), .A0N(cal_out[206]), .A1N(n5209), 
        .Y(n2205) );
  OAI2BB2X1 U9148 ( .B0(n5936), .B1(n5612), .A0N(cal_out[246]), .A1N(n5213), 
        .Y(n2165) );
  OAI2BB2X1 U9149 ( .B0(n5936), .B1(n5615), .A0N(cal_out[286]), .A1N(n5217), 
        .Y(n2125) );
  OAI2BB2X1 U9150 ( .B0(n5936), .B1(n5618), .A0N(cal_out[326]), .A1N(n5221), 
        .Y(n2085) );
  OAI2BB2X1 U9151 ( .B0(n5936), .B1(n5621), .A0N(cal_out[366]), .A1N(n5225), 
        .Y(n2045) );
  OAI2BB2X1 U9152 ( .B0(n5936), .B1(n5624), .A0N(cal_out[406]), .A1N(n5229), 
        .Y(n2005) );
  OAI2BB2X1 U9153 ( .B0(n5936), .B1(n5627), .A0N(cal_out[446]), .A1N(n5233), 
        .Y(n1965) );
  OAI2BB2X1 U9154 ( .B0(n5936), .B1(n5631), .A0N(cal_out[486]), .A1N(n5237), 
        .Y(n1925) );
  OAI2BB2X1 U9155 ( .B0(n5936), .B1(n5635), .A0N(cal_out[526]), .A1N(n5243), 
        .Y(n1885) );
  OAI2BB2X1 U9156 ( .B0(n5962), .B1(n5595), .A0N(cal_out[30]), .A1N(n5191), 
        .Y(n2381) );
  OAI2BB2X1 U9157 ( .B0(n5962), .B1(n5598), .A0N(cal_out[70]), .A1N(n5195), 
        .Y(n2341) );
  OAI2BB2X1 U9158 ( .B0(n5962), .B1(n5601), .A0N(cal_out[110]), .A1N(n5199), 
        .Y(n2301) );
  OAI2BB2X1 U9159 ( .B0(n5962), .B1(n5604), .A0N(cal_out[150]), .A1N(n5203), 
        .Y(n2261) );
  OAI2BB2X1 U9160 ( .B0(n5962), .B1(n5607), .A0N(cal_out[190]), .A1N(n5207), 
        .Y(n2221) );
  OAI2BB2X1 U9161 ( .B0(n5962), .B1(n5610), .A0N(cal_out[230]), .A1N(n5211), 
        .Y(n2181) );
  OAI2BB2X1 U9162 ( .B0(n5962), .B1(n5613), .A0N(cal_out[270]), .A1N(n5215), 
        .Y(n2141) );
  OAI2BB2X1 U9163 ( .B0(n5962), .B1(n5616), .A0N(cal_out[310]), .A1N(n5219), 
        .Y(n2101) );
  OAI2BB2X1 U9164 ( .B0(n5962), .B1(n5619), .A0N(cal_out[350]), .A1N(n5223), 
        .Y(n2061) );
  OAI2BB2X1 U9165 ( .B0(n5962), .B1(n5622), .A0N(cal_out[390]), .A1N(n5227), 
        .Y(n2021) );
  OAI2BB2X1 U9166 ( .B0(n5962), .B1(n5625), .A0N(cal_out[430]), .A1N(n5231), 
        .Y(n1981) );
  OAI2BB2X1 U9167 ( .B0(n5962), .B1(n5628), .A0N(cal_out[470]), .A1N(n5235), 
        .Y(n1941) );
  OAI2BB2X1 U9168 ( .B0(n5962), .B1(n5631), .A0N(cal_out[510]), .A1N(n5239), 
        .Y(n1901) );
  OAI2BB2X1 U9169 ( .B0(n5962), .B1(n5633), .A0N(cal_out[550]), .A1N(n5242), 
        .Y(n1861) );
  OAI2BB2X1 U9170 ( .B0(n5945), .B1(n5596), .A0N(cal_out[14]), .A1N(n5190), 
        .Y(n2397) );
  OAI2BB2X1 U9171 ( .B0(n5945), .B1(n5599), .A0N(cal_out[54]), .A1N(n5194), 
        .Y(n2357) );
  OAI2BB2X1 U9172 ( .B0(n5945), .B1(n5602), .A0N(cal_out[94]), .A1N(n5198), 
        .Y(n2317) );
  OAI2BB2X1 U9173 ( .B0(n5945), .B1(n5605), .A0N(cal_out[134]), .A1N(n5202), 
        .Y(n2277) );
  OAI2BB2X1 U9174 ( .B0(n5945), .B1(n5608), .A0N(cal_out[174]), .A1N(n5206), 
        .Y(n2237) );
  OAI2BB2X1 U9175 ( .B0(n5945), .B1(n5611), .A0N(cal_out[214]), .A1N(n5210), 
        .Y(n2197) );
  OAI2BB2X1 U9176 ( .B0(n5945), .B1(n5614), .A0N(cal_out[254]), .A1N(n5214), 
        .Y(n2157) );
  OAI2BB2X1 U9177 ( .B0(n5945), .B1(n5617), .A0N(cal_out[294]), .A1N(n5218), 
        .Y(n2117) );
  OAI2BB2X1 U9178 ( .B0(n5945), .B1(n5620), .A0N(cal_out[334]), .A1N(n5222), 
        .Y(n2077) );
  OAI2BB2X1 U9179 ( .B0(n5945), .B1(n5623), .A0N(cal_out[374]), .A1N(n5226), 
        .Y(n2037) );
  OAI2BB2X1 U9180 ( .B0(n5945), .B1(n5626), .A0N(cal_out[414]), .A1N(n5230), 
        .Y(n1997) );
  OAI2BB2X1 U9181 ( .B0(n5945), .B1(n5629), .A0N(cal_out[454]), .A1N(n5234), 
        .Y(n1957) );
  OAI2BB2X1 U9182 ( .B0(n5945), .B1(n5632), .A0N(cal_out[494]), .A1N(n5238), 
        .Y(n1917) );
  OAI2BB2X1 U9183 ( .B0(n5945), .B1(n5634), .A0N(cal_out[534]), .A1N(n5241), 
        .Y(n1877) );
  OAI2BB2X1 U9184 ( .B0(n5932), .B1(n5595), .A0N(cal_out[2]), .A1N(n5189), .Y(
        n2409) );
  OAI2BB2X1 U9185 ( .B0(n5932), .B1(n5598), .A0N(cal_out[42]), .A1N(n5193), 
        .Y(n2369) );
  OAI2BB2X1 U9186 ( .B0(n5932), .B1(n5601), .A0N(cal_out[82]), .A1N(n5197), 
        .Y(n2329) );
  OAI2BB2X1 U9187 ( .B0(n5932), .B1(n5604), .A0N(cal_out[122]), .A1N(n5201), 
        .Y(n2289) );
  OAI2BB2X1 U9188 ( .B0(n5932), .B1(n5607), .A0N(cal_out[162]), .A1N(n5205), 
        .Y(n2249) );
  OAI2BB2X1 U9189 ( .B0(n5932), .B1(n5610), .A0N(cal_out[202]), .A1N(n5209), 
        .Y(n2209) );
  OAI2BB2X1 U9190 ( .B0(n5932), .B1(n5613), .A0N(cal_out[242]), .A1N(n5213), 
        .Y(n2169) );
  OAI2BB2X1 U9191 ( .B0(n5932), .B1(n5616), .A0N(cal_out[282]), .A1N(n5217), 
        .Y(n2129) );
  OAI2BB2X1 U9192 ( .B0(n5932), .B1(n5619), .A0N(cal_out[322]), .A1N(n5221), 
        .Y(n2089) );
  OAI2BB2X1 U9193 ( .B0(n5932), .B1(n5622), .A0N(cal_out[362]), .A1N(n5225), 
        .Y(n2049) );
  OAI2BB2X1 U9194 ( .B0(n5932), .B1(n5625), .A0N(cal_out[402]), .A1N(n5229), 
        .Y(n2009) );
  OAI2BB2X1 U9195 ( .B0(n5932), .B1(n5628), .A0N(cal_out[442]), .A1N(n5233), 
        .Y(n1969) );
  OAI2BB2X1 U9196 ( .B0(n5932), .B1(n5631), .A0N(cal_out[482]), .A1N(n5237), 
        .Y(n1929) );
  OAI2BB2X1 U9197 ( .B0(n5932), .B1(n5635), .A0N(cal_out[522]), .A1N(n5243), 
        .Y(n1889) );
  OAI2BB2XL U9198 ( .B0(n5637), .B1(n5939), .A0N(cal_out[569]), .A1N(n5245), 
        .Y(n1842) );
  OAI2BB2XL U9199 ( .B0(n5636), .B1(n5950), .A0N(cal_out[579]), .A1N(n5246), 
        .Y(n1832) );
  OAI2BB2XL U9200 ( .B0(n5636), .B1(n5954), .A0N(cal_out[583]), .A1N(n5246), 
        .Y(n1828) );
  OAI2BB2XL U9201 ( .B0(n5636), .B1(n5951), .A0N(cal_out[580]), .A1N(n5246), 
        .Y(n1831) );
  OAI2BB2XL U9202 ( .B0(n5636), .B1(n5959), .A0N(cal_out[587]), .A1N(n5247), 
        .Y(n1824) );
  OAI2BB2XL U9203 ( .B0(n5636), .B1(n5960), .A0N(cal_out[588]), .A1N(n5247), 
        .Y(n1823) );
  OAI2BB2XL U9204 ( .B0(n5636), .B1(n5953), .A0N(cal_out[582]), .A1N(n5246), 
        .Y(n1829) );
  OAI2BB2XL U9205 ( .B0(n5637), .B1(n5935), .A0N(cal_out[565]), .A1N(n5245), 
        .Y(n1846) );
  OAI2BB2XL U9206 ( .B0(n5637), .B1(n5934), .A0N(cal_out[564]), .A1N(n5245), 
        .Y(n1847) );
  OAI2BB2XL U9207 ( .B0(n5636), .B1(n5957), .A0N(cal_out[585]), .A1N(n5247), 
        .Y(n1826) );
  OAI2BB2XL U9208 ( .B0(n5636), .B1(n5944), .A0N(cal_out[573]), .A1N(n5246), 
        .Y(n1838) );
  OAI2BB2XL U9209 ( .B0(n5637), .B1(n5938), .A0N(cal_out[568]), .A1N(n5245), 
        .Y(n1843) );
  OAI2BB2XL U9210 ( .B0(n5637), .B1(n5931), .A0N(cal_out[561]), .A1N(n5245), 
        .Y(n1850) );
  OAI2BB2XL U9211 ( .B0(n5636), .B1(n5961), .A0N(cal_out[589]), .A1N(n5247), 
        .Y(n1822) );
  OAI2BB2XL U9212 ( .B0(n5636), .B1(n5958), .A0N(cal_out[586]), .A1N(n5247), 
        .Y(n1825) );
  OAI2BB2XL U9213 ( .B0(n5636), .B1(n5955), .A0N(cal_out[584]), .A1N(n5247), 
        .Y(n1827) );
  OAI2BB2XL U9214 ( .B0(n5636), .B1(n5946), .A0N(cal_out[575]), .A1N(n5246), 
        .Y(n1836) );
  OAI2BB2XL U9215 ( .B0(n5637), .B1(n5942), .A0N(cal_out[571]), .A1N(n5245), 
        .Y(n1840) );
  OAI2BB2XL U9216 ( .B0(n5636), .B1(n5947), .A0N(cal_out[576]), .A1N(n5246), 
        .Y(n1835) );
  OAI2BB2XL U9217 ( .B0(n5637), .B1(n5940), .A0N(cal_out[570]), .A1N(n5245), 
        .Y(n1841) );
  OAI2BB2XL U9218 ( .B0(n5636), .B1(n5949), .A0N(cal_out[578]), .A1N(n5246), 
        .Y(n1833) );
  OAI2BB2XL U9219 ( .B0(n5637), .B1(n5937), .A0N(cal_out[567]), .A1N(n5245), 
        .Y(n1844) );
  OAI2BB2XL U9220 ( .B0(n5637), .B1(n5943), .A0N(cal_out[572]), .A1N(n5246), 
        .Y(n1839) );
  OAI2BB2XL U9221 ( .B0(n5636), .B1(n5930), .A0N(cal_out[560]), .A1N(n5245), 
        .Y(n1851) );
  OAI2BB2XL U9222 ( .B0(n5637), .B1(n5936), .A0N(cal_out[566]), .A1N(n5245), 
        .Y(n1845) );
  OAI2BB2XL U9223 ( .B0(n5637), .B1(n5962), .A0N(cal_out[590]), .A1N(n5247), 
        .Y(n1821) );
  OAI2BB2XL U9224 ( .B0(n5636), .B1(n5945), .A0N(cal_out[574]), .A1N(n5246), 
        .Y(n1837) );
  OAI2BB2XL U9225 ( .B0(n5637), .B1(n5932), .A0N(cal_out[562]), .A1N(n5245), 
        .Y(n1849) );
  NAND2X1 U9226 ( .A(c_plus[36]), .B(n779), .Y(n781) );
  NAND2X1 U9227 ( .A(c_plus[33]), .B(n828), .Y(n778) );
  NOR3X1 U9228 ( .A(cal_cnt[0]), .B(n5087), .C(n5892), .Y(n1516) );
  CLKINVX3 U9229 ( .A(n1013), .Y(n5861) );
  AOI22X1 U9230 ( .A0(n5052), .A1(in_addr_cnt[7]), .B0(calweight_addr[7]), 
        .B1(n5066), .Y(n1013) );
  CLKINVX3 U9231 ( .A(n1016), .Y(n5863) );
  AOI22X1 U9232 ( .A0(n5052), .A1(in_addr_cnt[5]), .B0(calweight_addr[5]), 
        .B1(n5066), .Y(n1016) );
  CLKINVX3 U9233 ( .A(n1022), .Y(n5869) );
  AOI22X1 U9234 ( .A0(n5052), .A1(in_addr_cnt[7]), .B0(calin_addr[7]), .B1(
        n5066), .Y(n1022) );
  CLKINVX3 U9235 ( .A(n1024), .Y(n5871) );
  AOI22X1 U9236 ( .A0(n5052), .A1(in_addr_cnt[5]), .B0(calin_addr[5]), .B1(
        n5066), .Y(n1024) );
  CLKINVX3 U9237 ( .A(n1019), .Y(n5866) );
  AOI22X1 U9238 ( .A0(n5051), .A1(in_addr_cnt[2]), .B0(calweight_addr[2]), 
        .B1(n5066), .Y(n1019) );
  CLKINVX3 U9239 ( .A(n1027), .Y(n5874) );
  AOI22X1 U9240 ( .A0(n5051), .A1(in_addr_cnt[2]), .B0(calin_addr[2]), .B1(
        n5066), .Y(n1027) );
  CMPR22X1 U9241 ( .A(in_cnt_64[1]), .B(in_cnt_64[0]), .CO(add_220_carry[2]), 
        .S(N1035) );
  CLKINVX3 U9242 ( .A(n1018), .Y(n5865) );
  AOI22X1 U9243 ( .A0(n5052), .A1(in_addr_cnt[3]), .B0(calweight_addr[3]), 
        .B1(n5066), .Y(n1018) );
  CLKINVX3 U9244 ( .A(n1026), .Y(n5873) );
  AOI22X1 U9245 ( .A0(n5052), .A1(in_addr_cnt[3]), .B0(calin_addr[3]), .B1(
        n5066), .Y(n1026) );
  CLKINVX3 U9246 ( .A(n1020), .Y(n5867) );
  AOI22X1 U9247 ( .A0(n5052), .A1(in_addr_cnt[1]), .B0(calweight_addr[1]), 
        .B1(n5066), .Y(n1020) );
  CLKINVX3 U9248 ( .A(n1028), .Y(n5875) );
  AOI22X1 U9249 ( .A0(n5052), .A1(in_addr_cnt[1]), .B0(calin_addr[1]), .B1(
        n5066), .Y(n1028) );
  OAI2BB2X1 U9250 ( .B0(n5594), .B1(n5970), .A0N(cal_out[39]), .A1N(n5190), 
        .Y(n2372) );
  OAI2BB2X1 U9251 ( .B0(n5597), .B1(n5970), .A0N(cal_out[79]), .A1N(n5194), 
        .Y(n2332) );
  OAI2BB2X1 U9252 ( .B0(n5600), .B1(n5970), .A0N(cal_out[119]), .A1N(n5198), 
        .Y(n2292) );
  OAI2BB2X1 U9253 ( .B0(n5603), .B1(n5970), .A0N(cal_out[159]), .A1N(n5202), 
        .Y(n2252) );
  OAI2BB2X1 U9254 ( .B0(n5606), .B1(n5970), .A0N(cal_out[199]), .A1N(n5206), 
        .Y(n2212) );
  OAI2BB2X1 U9255 ( .B0(n5609), .B1(n5970), .A0N(cal_out[239]), .A1N(n5210), 
        .Y(n2172) );
  OAI2BB2X1 U9256 ( .B0(n5612), .B1(n5970), .A0N(cal_out[279]), .A1N(n5214), 
        .Y(n2132) );
  OAI2BB2X1 U9257 ( .B0(n5615), .B1(n5970), .A0N(cal_out[319]), .A1N(n5218), 
        .Y(n2092) );
  OAI2BB2X1 U9258 ( .B0(n5618), .B1(n5970), .A0N(cal_out[359]), .A1N(n5222), 
        .Y(n2052) );
  OAI2BB2X1 U9259 ( .B0(n5621), .B1(n5970), .A0N(cal_out[399]), .A1N(n5226), 
        .Y(n2012) );
  OAI2BB2X1 U9260 ( .B0(n5624), .B1(n5970), .A0N(cal_out[439]), .A1N(n5230), 
        .Y(n1972) );
  OAI2BB2X1 U9261 ( .B0(n5627), .B1(n5970), .A0N(cal_out[479]), .A1N(n5235), 
        .Y(n1932) );
  OAI2BB2X1 U9262 ( .B0(n5630), .B1(n5970), .A0N(cal_out[519]), .A1N(n5238), 
        .Y(n1892) );
  OAI2BB2X1 U9263 ( .B0(n5633), .B1(n5970), .A0N(cal_out[559]), .A1N(n5243), 
        .Y(n1852) );
  OAI2BB2X1 U9264 ( .B0(n757), .B1(n5970), .A0N(cal_out[599]), .A1N(n5857), 
        .Y(n1812) );
  CMPR22X1 U9265 ( .A(in_cnt_64[2]), .B(add_220_carry[2]), .CO(
        add_220_carry[3]), .S(N1036) );
  CMPR22X1 U9266 ( .A(in_cnt_64[3]), .B(add_220_carry[3]), .CO(
        add_220_carry[4]), .S(N1037) );
  OAI2BB2X1 U9267 ( .B0(n5594), .B1(n5085), .A0N(cal_out[31]), .A1N(n5191), 
        .Y(n2380) );
  OAI2BB2X1 U9268 ( .B0(n5597), .B1(n5085), .A0N(cal_out[71]), .A1N(n5195), 
        .Y(n2340) );
  OAI2BB2X1 U9269 ( .B0(n5600), .B1(n5085), .A0N(cal_out[111]), .A1N(n5199), 
        .Y(n2300) );
  OAI2BB2X1 U9270 ( .B0(n5603), .B1(n5085), .A0N(cal_out[151]), .A1N(n5203), 
        .Y(n2260) );
  OAI2BB2X1 U9271 ( .B0(n5606), .B1(n5085), .A0N(cal_out[191]), .A1N(n5207), 
        .Y(n2220) );
  OAI2BB2X1 U9272 ( .B0(n5609), .B1(n5085), .A0N(cal_out[231]), .A1N(n5211), 
        .Y(n2180) );
  OAI2BB2X1 U9273 ( .B0(n5612), .B1(n5085), .A0N(cal_out[271]), .A1N(n5215), 
        .Y(n2140) );
  OAI2BB2X1 U9274 ( .B0(n5615), .B1(n5085), .A0N(cal_out[311]), .A1N(n5219), 
        .Y(n2100) );
  OAI2BB2X1 U9275 ( .B0(n5618), .B1(n5085), .A0N(cal_out[351]), .A1N(n5223), 
        .Y(n2060) );
  OAI2BB2X1 U9276 ( .B0(n5621), .B1(n5085), .A0N(cal_out[391]), .A1N(n5227), 
        .Y(n2020) );
  OAI2BB2X1 U9277 ( .B0(n5624), .B1(n5085), .A0N(cal_out[431]), .A1N(n5231), 
        .Y(n1980) );
  OAI2BB2X1 U9278 ( .B0(n5627), .B1(n5085), .A0N(cal_out[471]), .A1N(n5235), 
        .Y(n1940) );
  OAI2BB2X1 U9279 ( .B0(n5630), .B1(n5085), .A0N(cal_out[511]), .A1N(n5239), 
        .Y(n1900) );
  OAI2BB2X1 U9280 ( .B0(n5633), .B1(n5085), .A0N(cal_out[551]), .A1N(n5242), 
        .Y(n1860) );
  OAI2BB2X1 U9281 ( .B0(n5637), .B1(n5085), .A0N(cal_out[591]), .A1N(n5247), 
        .Y(n1820) );
  OAI2BB2X1 U9282 ( .B0(n757), .B1(n5966), .A0N(cal_out[595]), .A1N(n5247), 
        .Y(n1816) );
  OAI2BB2X1 U9283 ( .B0(n5636), .B1(n5952), .A0N(cal_out[581]), .A1N(n5246), 
        .Y(n1830) );
  OAI2BB2X1 U9284 ( .B0(n5933), .B1(n5596), .A0N(cal_out[3]), .A1N(n5189), .Y(
        n2408) );
  OAI2BB2X1 U9285 ( .B0(n5933), .B1(n5599), .A0N(cal_out[43]), .A1N(n5193), 
        .Y(n2368) );
  OAI2BB2X1 U9286 ( .B0(n5933), .B1(n5602), .A0N(cal_out[83]), .A1N(n5197), 
        .Y(n2328) );
  OAI2BB2X1 U9287 ( .B0(n5933), .B1(n5605), .A0N(cal_out[123]), .A1N(n5201), 
        .Y(n2288) );
  OAI2BB2X1 U9288 ( .B0(n5933), .B1(n5608), .A0N(cal_out[163]), .A1N(n5205), 
        .Y(n2248) );
  OAI2BB2X1 U9289 ( .B0(n5933), .B1(n5611), .A0N(cal_out[203]), .A1N(n5209), 
        .Y(n2208) );
  OAI2BB2X1 U9290 ( .B0(n5933), .B1(n5614), .A0N(cal_out[243]), .A1N(n5213), 
        .Y(n2168) );
  OAI2BB2X1 U9291 ( .B0(n5933), .B1(n5617), .A0N(cal_out[283]), .A1N(n5217), 
        .Y(n2128) );
  OAI2BB2X1 U9292 ( .B0(n5933), .B1(n5620), .A0N(cal_out[323]), .A1N(n5221), 
        .Y(n2088) );
  OAI2BB2X1 U9293 ( .B0(n5933), .B1(n5623), .A0N(cal_out[363]), .A1N(n5225), 
        .Y(n2048) );
  OAI2BB2X1 U9294 ( .B0(n5933), .B1(n5626), .A0N(cal_out[403]), .A1N(n5229), 
        .Y(n2008) );
  OAI2BB2X1 U9295 ( .B0(n5933), .B1(n5629), .A0N(cal_out[443]), .A1N(n5233), 
        .Y(n1968) );
  OAI2BB2X1 U9296 ( .B0(n5933), .B1(n5632), .A0N(cal_out[483]), .A1N(n5237), 
        .Y(n1928) );
  OAI2BB2X1 U9297 ( .B0(n5933), .B1(n5635), .A0N(cal_out[523]), .A1N(n5241), 
        .Y(n1888) );
  OAI2BB2X1 U9298 ( .B0(n5637), .B1(n5933), .A0N(cal_out[563]), .A1N(n5245), 
        .Y(n1848) );
  OAI2BB2X1 U9299 ( .B0(n5966), .B1(n5595), .A0N(cal_out[35]), .A1N(n5191), 
        .Y(n2376) );
  OAI2BB2X1 U9300 ( .B0(n5966), .B1(n5598), .A0N(cal_out[75]), .A1N(n5195), 
        .Y(n2336) );
  OAI2BB2X1 U9301 ( .B0(n5966), .B1(n5601), .A0N(cal_out[115]), .A1N(n5199), 
        .Y(n2296) );
  OAI2BB2X1 U9302 ( .B0(n5966), .B1(n5604), .A0N(cal_out[155]), .A1N(n5203), 
        .Y(n2256) );
  OAI2BB2X1 U9303 ( .B0(n5966), .B1(n5607), .A0N(cal_out[195]), .A1N(n5207), 
        .Y(n2216) );
  OAI2BB2X1 U9304 ( .B0(n5966), .B1(n5610), .A0N(cal_out[235]), .A1N(n5211), 
        .Y(n2176) );
  OAI2BB2X1 U9305 ( .B0(n5966), .B1(n5613), .A0N(cal_out[275]), .A1N(n5215), 
        .Y(n2136) );
  OAI2BB2X1 U9306 ( .B0(n5966), .B1(n5616), .A0N(cal_out[315]), .A1N(n5219), 
        .Y(n2096) );
  OAI2BB2X1 U9307 ( .B0(n5966), .B1(n5619), .A0N(cal_out[355]), .A1N(n5223), 
        .Y(n2056) );
  OAI2BB2X1 U9308 ( .B0(n5966), .B1(n5622), .A0N(cal_out[395]), .A1N(n5227), 
        .Y(n2016) );
  OAI2BB2X1 U9309 ( .B0(n5966), .B1(n5625), .A0N(cal_out[435]), .A1N(n5231), 
        .Y(n1976) );
  OAI2BB2X1 U9310 ( .B0(n5966), .B1(n5628), .A0N(cal_out[475]), .A1N(n5235), 
        .Y(n1936) );
  OAI2BB2X1 U9311 ( .B0(n5966), .B1(n5631), .A0N(cal_out[515]), .A1N(n5239), 
        .Y(n1896) );
  OAI2BB2X1 U9312 ( .B0(n5966), .B1(n5634), .A0N(cal_out[555]), .A1N(n5242), 
        .Y(n1856) );
  OAI2BB2X1 U9313 ( .B0(n5636), .B1(n5948), .A0N(cal_out[577]), .A1N(n5246), 
        .Y(n1834) );
  OAI2BB2X1 U9314 ( .B0(n5964), .B1(n5594), .A0N(cal_out[33]), .A1N(n5191), 
        .Y(n2378) );
  OAI2BB2X1 U9315 ( .B0(n5964), .B1(n5597), .A0N(cal_out[73]), .A1N(n5195), 
        .Y(n2338) );
  OAI2BB2X1 U9316 ( .B0(n5964), .B1(n5600), .A0N(cal_out[113]), .A1N(n5199), 
        .Y(n2298) );
  OAI2BB2X1 U9317 ( .B0(n5964), .B1(n5603), .A0N(cal_out[153]), .A1N(n5203), 
        .Y(n2258) );
  OAI2BB2X1 U9318 ( .B0(n5964), .B1(n5606), .A0N(cal_out[193]), .A1N(n5207), 
        .Y(n2218) );
  OAI2BB2X1 U9319 ( .B0(n5964), .B1(n5609), .A0N(cal_out[233]), .A1N(n5211), 
        .Y(n2178) );
  OAI2BB2X1 U9320 ( .B0(n5964), .B1(n5612), .A0N(cal_out[273]), .A1N(n5215), 
        .Y(n2138) );
  OAI2BB2X1 U9321 ( .B0(n5964), .B1(n5615), .A0N(cal_out[313]), .A1N(n5219), 
        .Y(n2098) );
  OAI2BB2X1 U9322 ( .B0(n5964), .B1(n5618), .A0N(cal_out[353]), .A1N(n5223), 
        .Y(n2058) );
  OAI2BB2X1 U9323 ( .B0(n5964), .B1(n5621), .A0N(cal_out[393]), .A1N(n5227), 
        .Y(n2018) );
  OAI2BB2X1 U9324 ( .B0(n5964), .B1(n5624), .A0N(cal_out[433]), .A1N(n5231), 
        .Y(n1978) );
  OAI2BB2X1 U9325 ( .B0(n5964), .B1(n5627), .A0N(cal_out[473]), .A1N(n5235), 
        .Y(n1938) );
  OAI2BB2X1 U9326 ( .B0(n5964), .B1(n5630), .A0N(cal_out[513]), .A1N(n5239), 
        .Y(n1898) );
  OAI2BB2X1 U9327 ( .B0(n5964), .B1(n5633), .A0N(cal_out[553]), .A1N(n5242), 
        .Y(n1858) );
  OAI2BB2X1 U9328 ( .B0(n5964), .B1(n5636), .A0N(cal_out[593]), .A1N(n5247), 
        .Y(n1818) );
  OAI2BB2X1 U9329 ( .B0(n5952), .B1(n5595), .A0N(cal_out[21]), .A1N(n5190), 
        .Y(n2390) );
  OAI2BB2X1 U9330 ( .B0(n5952), .B1(n5598), .A0N(cal_out[61]), .A1N(n5194), 
        .Y(n2350) );
  OAI2BB2X1 U9331 ( .B0(n5952), .B1(n5601), .A0N(cal_out[101]), .A1N(n5198), 
        .Y(n2310) );
  OAI2BB2X1 U9332 ( .B0(n5952), .B1(n5604), .A0N(cal_out[141]), .A1N(n5202), 
        .Y(n2270) );
  OAI2BB2X1 U9333 ( .B0(n5952), .B1(n5607), .A0N(cal_out[181]), .A1N(n5206), 
        .Y(n2230) );
  OAI2BB2X1 U9334 ( .B0(n5952), .B1(n5610), .A0N(cal_out[221]), .A1N(n5210), 
        .Y(n2190) );
  OAI2BB2X1 U9335 ( .B0(n5952), .B1(n5613), .A0N(cal_out[261]), .A1N(n5214), 
        .Y(n2150) );
  OAI2BB2X1 U9336 ( .B0(n5952), .B1(n5616), .A0N(cal_out[301]), .A1N(n5218), 
        .Y(n2110) );
  OAI2BB2X1 U9337 ( .B0(n5952), .B1(n5619), .A0N(cal_out[341]), .A1N(n5222), 
        .Y(n2070) );
  OAI2BB2X1 U9338 ( .B0(n5952), .B1(n5622), .A0N(cal_out[381]), .A1N(n5226), 
        .Y(n2030) );
  OAI2BB2X1 U9339 ( .B0(n5952), .B1(n5625), .A0N(cal_out[421]), .A1N(n5230), 
        .Y(n1990) );
  OAI2BB2X1 U9340 ( .B0(n5952), .B1(n5628), .A0N(cal_out[461]), .A1N(n5234), 
        .Y(n1950) );
  OAI2BB2X1 U9341 ( .B0(n5952), .B1(n5631), .A0N(cal_out[501]), .A1N(n5238), 
        .Y(n1910) );
  OAI2BB2X1 U9342 ( .B0(n5952), .B1(n5634), .A0N(cal_out[541]), .A1N(n5241), 
        .Y(n1870) );
  OAI2BB2X1 U9343 ( .B0(n5084), .B1(n5637), .A0N(length_reg[89]), .A1N(n5857), 
        .Y(n1722) );
  OAI2BB2X1 U9344 ( .B0(n5948), .B1(n5596), .A0N(cal_out[17]), .A1N(n5190), 
        .Y(n2394) );
  OAI2BB2X1 U9345 ( .B0(n5948), .B1(n5599), .A0N(cal_out[57]), .A1N(n5194), 
        .Y(n2354) );
  OAI2BB2X1 U9346 ( .B0(n5948), .B1(n5602), .A0N(cal_out[97]), .A1N(n5198), 
        .Y(n2314) );
  OAI2BB2X1 U9347 ( .B0(n5948), .B1(n5605), .A0N(cal_out[137]), .A1N(n5202), 
        .Y(n2274) );
  OAI2BB2X1 U9348 ( .B0(n5948), .B1(n5608), .A0N(cal_out[177]), .A1N(n5206), 
        .Y(n2234) );
  OAI2BB2X1 U9349 ( .B0(n5948), .B1(n5611), .A0N(cal_out[217]), .A1N(n5210), 
        .Y(n2194) );
  OAI2BB2X1 U9350 ( .B0(n5948), .B1(n5614), .A0N(cal_out[257]), .A1N(n5214), 
        .Y(n2154) );
  OAI2BB2X1 U9351 ( .B0(n5948), .B1(n5617), .A0N(cal_out[297]), .A1N(n5218), 
        .Y(n2114) );
  OAI2BB2X1 U9352 ( .B0(n5948), .B1(n5620), .A0N(cal_out[337]), .A1N(n5222), 
        .Y(n2074) );
  OAI2BB2X1 U9353 ( .B0(n5948), .B1(n5623), .A0N(cal_out[377]), .A1N(n5226), 
        .Y(n2034) );
  OAI2BB2X1 U9354 ( .B0(n5948), .B1(n5626), .A0N(cal_out[417]), .A1N(n5230), 
        .Y(n1994) );
  OAI2BB2X1 U9355 ( .B0(n5948), .B1(n5629), .A0N(cal_out[457]), .A1N(n5234), 
        .Y(n1954) );
  OAI2BB2X1 U9356 ( .B0(n5948), .B1(n5632), .A0N(cal_out[497]), .A1N(n5238), 
        .Y(n1914) );
  OAI2BB2X1 U9357 ( .B0(n5948), .B1(n5634), .A0N(cal_out[537]), .A1N(n5241), 
        .Y(n1874) );
  OAI2BB2X1 U9358 ( .B0(n5084), .B1(n5595), .A0N(length_reg[5]), .A1N(n5189), 
        .Y(n1806) );
  OAI2BB2X1 U9359 ( .B0(n5084), .B1(n5598), .A0N(length_reg[11]), .A1N(n5193), 
        .Y(n1800) );
  OAI2BB2X1 U9360 ( .B0(n5084), .B1(n5601), .A0N(length_reg[17]), .A1N(n5197), 
        .Y(n1794) );
  OAI2BB2X1 U9361 ( .B0(n5084), .B1(n5604), .A0N(length_reg[23]), .A1N(n5201), 
        .Y(n1788) );
  OAI2BB2X1 U9362 ( .B0(n5084), .B1(n5607), .A0N(length_reg[29]), .A1N(n5205), 
        .Y(n1782) );
  OAI2BB2X1 U9363 ( .B0(n5084), .B1(n5610), .A0N(length_reg[35]), .A1N(n5209), 
        .Y(n1776) );
  OAI2BB2X1 U9364 ( .B0(n5084), .B1(n5613), .A0N(length_reg[41]), .A1N(n5213), 
        .Y(n1770) );
  OAI2BB2X1 U9365 ( .B0(n5084), .B1(n5616), .A0N(length_reg[47]), .A1N(n5217), 
        .Y(n1764) );
  OAI2BB2X1 U9366 ( .B0(n5084), .B1(n5619), .A0N(length_reg[53]), .A1N(n5221), 
        .Y(n1758) );
  OAI2BB2X1 U9367 ( .B0(n5084), .B1(n5622), .A0N(length_reg[59]), .A1N(n5225), 
        .Y(n1752) );
  OAI2BB2X1 U9368 ( .B0(n5084), .B1(n5625), .A0N(length_reg[65]), .A1N(n5229), 
        .Y(n1746) );
  OAI2BB2X1 U9369 ( .B0(n5084), .B1(n5628), .A0N(length_reg[71]), .A1N(n5234), 
        .Y(n1740) );
  OAI2BB2X1 U9370 ( .B0(n5084), .B1(n5631), .A0N(length_reg[77]), .A1N(n5237), 
        .Y(n1734) );
  OAI2BB2X1 U9371 ( .B0(n5084), .B1(n5633), .A0N(length_reg[83]), .A1N(n5243), 
        .Y(n1728) );
  OAI2BB2X1 U9372 ( .B0(n757), .B1(n5968), .A0N(cal_out[597]), .A1N(n5857), 
        .Y(n1814) );
  OAI2BB2X1 U9373 ( .B0(n757), .B1(n5969), .A0N(cal_out[598]), .A1N(n5857), 
        .Y(n1813) );
  OAI2BB2X1 U9374 ( .B0(n5969), .B1(n5594), .A0N(cal_out[38]), .A1N(n5843), 
        .Y(n2373) );
  OAI2BB2X1 U9375 ( .B0(n5969), .B1(n5597), .A0N(cal_out[78]), .A1N(n5844), 
        .Y(n2333) );
  OAI2BB2X1 U9376 ( .B0(n5969), .B1(n5600), .A0N(cal_out[118]), .A1N(n5845), 
        .Y(n2293) );
  OAI2BB2X1 U9377 ( .B0(n5969), .B1(n5603), .A0N(cal_out[158]), .A1N(n5846), 
        .Y(n2253) );
  OAI2BB2X1 U9378 ( .B0(n5969), .B1(n5606), .A0N(cal_out[198]), .A1N(n5847), 
        .Y(n2213) );
  OAI2BB2X1 U9379 ( .B0(n5969), .B1(n5609), .A0N(cal_out[238]), .A1N(n5848), 
        .Y(n2173) );
  OAI2BB2X1 U9380 ( .B0(n5969), .B1(n5612), .A0N(cal_out[278]), .A1N(n5849), 
        .Y(n2133) );
  OAI2BB2X1 U9381 ( .B0(n5969), .B1(n5615), .A0N(cal_out[318]), .A1N(n5850), 
        .Y(n2093) );
  OAI2BB2X1 U9382 ( .B0(n5969), .B1(n5618), .A0N(cal_out[358]), .A1N(n5851), 
        .Y(n2053) );
  OAI2BB2X1 U9383 ( .B0(n5969), .B1(n5621), .A0N(cal_out[398]), .A1N(n5852), 
        .Y(n2013) );
  OAI2BB2X1 U9384 ( .B0(n5969), .B1(n5624), .A0N(cal_out[438]), .A1N(n5853), 
        .Y(n1973) );
  OAI2BB2X1 U9385 ( .B0(n5969), .B1(n5627), .A0N(cal_out[478]), .A1N(n5854), 
        .Y(n1933) );
  OAI2BB2X1 U9386 ( .B0(n5969), .B1(n5630), .A0N(cal_out[518]), .A1N(n5855), 
        .Y(n1893) );
  OAI2BB2X1 U9387 ( .B0(n5969), .B1(n5633), .A0N(cal_out[558]), .A1N(n5243), 
        .Y(n1853) );
  OAI2BB2X1 U9388 ( .B0(n5968), .B1(n5594), .A0N(cal_out[37]), .A1N(n5843), 
        .Y(n2374) );
  OAI2BB2X1 U9389 ( .B0(n5968), .B1(n5597), .A0N(cal_out[77]), .A1N(n5844), 
        .Y(n2334) );
  OAI2BB2X1 U9390 ( .B0(n5968), .B1(n5600), .A0N(cal_out[117]), .A1N(n5845), 
        .Y(n2294) );
  OAI2BB2X1 U9391 ( .B0(n5968), .B1(n5603), .A0N(cal_out[157]), .A1N(n5846), 
        .Y(n2254) );
  OAI2BB2X1 U9392 ( .B0(n5968), .B1(n5606), .A0N(cal_out[197]), .A1N(n5847), 
        .Y(n2214) );
  OAI2BB2X1 U9393 ( .B0(n5968), .B1(n5609), .A0N(cal_out[237]), .A1N(n5848), 
        .Y(n2174) );
  OAI2BB2X1 U9394 ( .B0(n5968), .B1(n5612), .A0N(cal_out[277]), .A1N(n5849), 
        .Y(n2134) );
  OAI2BB2X1 U9395 ( .B0(n5968), .B1(n5615), .A0N(cal_out[317]), .A1N(n5850), 
        .Y(n2094) );
  OAI2BB2X1 U9396 ( .B0(n5968), .B1(n5618), .A0N(cal_out[357]), .A1N(n5851), 
        .Y(n2054) );
  OAI2BB2X1 U9397 ( .B0(n5968), .B1(n5621), .A0N(cal_out[397]), .A1N(n5852), 
        .Y(n2014) );
  OAI2BB2X1 U9398 ( .B0(n5968), .B1(n5624), .A0N(cal_out[437]), .A1N(n5853), 
        .Y(n1974) );
  OAI2BB2X1 U9399 ( .B0(n5968), .B1(n5627), .A0N(cal_out[477]), .A1N(n5854), 
        .Y(n1934) );
  OAI2BB2X1 U9400 ( .B0(n5968), .B1(n5630), .A0N(cal_out[517]), .A1N(n5855), 
        .Y(n1894) );
  OAI2BB2X1 U9401 ( .B0(n5968), .B1(n5633), .A0N(cal_out[557]), .A1N(n5243), 
        .Y(n1854) );
  NAND2X1 U9402 ( .A(m_size[0]), .B(m_size[1]), .Y(calout_num_0_) );
  OAI21XL U9403 ( .A0(n744), .A1(n5978), .B0(n745), .Y(n1718) );
  AOI21X1 U9404 ( .A0(n5878), .A1(n4889), .B0(n742), .Y(n744) );
  NAND4X1 U9405 ( .A(n741), .B(N944), .C(N943), .D(n5978), .Y(n745) );
  INVX1 U9406 ( .A(N945), .Y(n5978) );
  XNOR2X1 U9407 ( .A(in_addr_cnt[7]), .B(N1233), .Y(n983) );
  INVX1 U9408 ( .A(n740), .Y(n5840) );
  AOI32X1 U9409 ( .A0(n741), .A1(n4889), .A2(N943), .B0(n742), .B1(N944), .Y(
        n740) );
  AND2X2 U9410 ( .A(N1361), .B(n5250), .Y(N1369) );
  XNOR2X1 U9411 ( .A(in_addr_cnt[5]), .B(n5662), .Y(n985) );
  NAND2BX1 U9412 ( .AN(n752), .B(n750), .Y(n1721) );
  OAI32X1 U9413 ( .A0(n727), .A1(out_cnt_6[2]), .A2(n748), .B0(n726), .B1(n749), .Y(n752) );
  XNOR2X1 U9414 ( .A(out_cnt_6[2]), .B(N14321), .Y(n1089) );
  XNOR2XL U9415 ( .A(in_addr_cnt[4]), .B(n5662), .Y(n989) );
  NOR2X1 U9416 ( .A(N14321), .B(n1089), .Y(n1088) );
  NAND2X1 U9417 ( .A(n751), .B(n750), .Y(n1720) );
  XNOR2X1 U9418 ( .A(n5972), .B(out_cnt_6[0]), .Y(n751) );
  NAND2X1 U9419 ( .A(n5972), .B(out_cnt_6[0]), .Y(n748) );
  OAI32X1 U9420 ( .A0(n746), .A1(N942), .A2(n747), .B0(n4890), .B1(n5879), .Y(
        n4472) );
  INVX1 U9421 ( .A(n747), .Y(n5879) );
  BUFX3 U9422 ( .A(cal_cnt[3]), .Y(n5086) );
  OAI2BB1X1 U9423 ( .A0N(N12206), .A1N(n5062), .B0(n1178), .Y(N12566) );
  AOI22X1 U9424 ( .A0(N12086), .A1(n1138), .B0(N12486), .B1(n1139), .Y(n1178)
         );
  AND4X2 U9425 ( .A(n843), .B(n844), .C(n845), .D(n846), .Y(n803) );
  NOR3X1 U9426 ( .A(n849), .B(c_plus[23]), .C(c_plus[13]), .Y(n844) );
  NOR3X1 U9427 ( .A(n847), .B(c_plus[34]), .C(c_plus[33]), .Y(n846) );
  NOR3X1 U9428 ( .A(n848), .B(c_plus[28]), .C(c_plus[27]), .Y(n845) );
  OAI221XL U9429 ( .A0(N14321), .A1(n748), .B0(n749), .B1(n727), .C0(n750), 
        .Y(n1719) );
  ADDHXL U9430 ( .A(in_cnt_64[4]), .B(add_220_carry[4]), .CO(add_220_carry[5]), 
        .S(N1038) );
  AND2X2 U9431 ( .A(N1354), .B(n5250), .Y(N1362) );
  NOR2X1 U9432 ( .A(n755), .B(n728), .Y(n749) );
  CMPR22X1 U9433 ( .A(in_matrix_cnt[1]), .B(in_matrix_cnt[0]), .CO(
        add_250_carry[2]), .S(N1086) );
  CMPR22X1 U9434 ( .A(in_matrix_cnt[2]), .B(add_250_carry[2]), .CO(
        add_250_carry[3]), .S(N1087) );
  NOR2X1 U9435 ( .A(N944), .B(N945), .Y(n4498) );
  NOR2X1 U9436 ( .A(n4489), .B(N942), .Y(n4506) );
  NOR2X1 U9437 ( .A(n4889), .B(N945), .Y(n4507) );
  NOR2X1 U9438 ( .A(n4890), .B(n4489), .Y(n4509) );
  AOI22X1 U9439 ( .A0(cal_out[519]), .A1(n4894), .B0(cal_out[319]), .B1(n4866), 
        .Y(n4503) );
  NOR2X1 U9440 ( .A(N942), .B(N943), .Y(n4504) );
  NOR2X1 U9441 ( .A(n4890), .B(N943), .Y(n4505) );
  AOI22X1 U9442 ( .A0(cal_out[599]), .A1(n4898), .B0(cal_out[559]), .B1(n4868), 
        .Y(n4502) );
  AND2X1 U9443 ( .A(N945), .B(N944), .Y(n4499) );
  AOI22X1 U9444 ( .A0(cal_out[39]), .A1(n4902), .B0(cal_out[479]), .B1(n4870), 
        .Y(n4501) );
  AOI22X1 U9445 ( .A0(cal_out[119]), .A1(n4906), .B0(cal_out[79]), .B1(n4872), 
        .Y(n4500) );
  NAND4X1 U9446 ( .A(n4503), .B(n4502), .C(n4501), .D(n4500), .Y(n4513) );
  AOI22X1 U9447 ( .A0(cal_out[439]), .A1(n4910), .B0(cal_out[399]), .B1(n4878), 
        .Y(n4512) );
  AND2X1 U9448 ( .A(N945), .B(n4889), .Y(n4508) );
  AND2X1 U9449 ( .A(n4508), .B(n4506), .Y(n4882) );
  AOI222X1 U9450 ( .A0(cal_out[199]), .A1(n4917), .B0(cal_out[279]), .B1(n4881), .C0(cal_out[239]), .C1(n4880), .Y(n4511) );
  AOI22X1 U9451 ( .A0(cal_out[359]), .A1(n4921), .B0(cal_out[159]), .B1(n4883), 
        .Y(n4510) );
  NAND4BXL U9452 ( .AN(n4513), .B(n4512), .C(n4511), .D(n4510), .Y(
        value_out[39]) );
  AOI22X1 U9453 ( .A0(cal_out[518]), .A1(n4894), .B0(cal_out[318]), .B1(n4866), 
        .Y(n4517) );
  AOI22X1 U9454 ( .A0(cal_out[598]), .A1(n4898), .B0(cal_out[558]), .B1(n4868), 
        .Y(n4516) );
  AOI22X1 U9455 ( .A0(cal_out[38]), .A1(n4902), .B0(cal_out[478]), .B1(n4870), 
        .Y(n4515) );
  AOI22X1 U9456 ( .A0(cal_out[118]), .A1(n4906), .B0(cal_out[78]), .B1(n4872), 
        .Y(n4514) );
  NAND4X1 U9457 ( .A(n4517), .B(n4516), .C(n4515), .D(n4514), .Y(n4521) );
  AOI22X1 U9458 ( .A0(cal_out[438]), .A1(n4910), .B0(cal_out[398]), .B1(n4878), 
        .Y(n4520) );
  AOI222X1 U9459 ( .A0(cal_out[198]), .A1(n4917), .B0(cal_out[278]), .B1(n4881), .C0(cal_out[238]), .C1(n4880), .Y(n4519) );
  AOI22X1 U9460 ( .A0(cal_out[358]), .A1(n4921), .B0(cal_out[158]), .B1(n4883), 
        .Y(n4518) );
  NAND4BXL U9461 ( .AN(n4521), .B(n4520), .C(n4519), .D(n4518), .Y(
        value_out[38]) );
  AOI22X1 U9462 ( .A0(cal_out[517]), .A1(n4894), .B0(cal_out[317]), .B1(n4866), 
        .Y(n4525) );
  AOI22X1 U9463 ( .A0(cal_out[597]), .A1(n4898), .B0(cal_out[557]), .B1(n4868), 
        .Y(n4524) );
  AOI22X1 U9464 ( .A0(cal_out[37]), .A1(n4902), .B0(cal_out[477]), .B1(n4870), 
        .Y(n4523) );
  AOI22X1 U9465 ( .A0(cal_out[117]), .A1(n4906), .B0(cal_out[77]), .B1(n4872), 
        .Y(n4522) );
  NAND4X1 U9466 ( .A(n4525), .B(n4524), .C(n4523), .D(n4522), .Y(n4529) );
  AOI22X1 U9467 ( .A0(cal_out[437]), .A1(n4910), .B0(cal_out[397]), .B1(n4878), 
        .Y(n4528) );
  AOI222X1 U9468 ( .A0(cal_out[197]), .A1(n4917), .B0(cal_out[277]), .B1(n4881), .C0(cal_out[237]), .C1(n4880), .Y(n4527) );
  AOI22X1 U9469 ( .A0(cal_out[357]), .A1(n4921), .B0(cal_out[157]), .B1(n4883), 
        .Y(n4526) );
  NAND4BXL U9470 ( .AN(n4529), .B(n4528), .C(n4527), .D(n4526), .Y(
        value_out[37]) );
  AOI22X1 U9471 ( .A0(cal_out[516]), .A1(n4894), .B0(cal_out[316]), .B1(n4866), 
        .Y(n4533) );
  AOI22X1 U9472 ( .A0(cal_out[596]), .A1(n4898), .B0(cal_out[556]), .B1(n4868), 
        .Y(n4532) );
  AOI22X1 U9473 ( .A0(cal_out[36]), .A1(n4902), .B0(cal_out[476]), .B1(n4870), 
        .Y(n4531) );
  AOI22X1 U9474 ( .A0(cal_out[116]), .A1(n4906), .B0(cal_out[76]), .B1(n4872), 
        .Y(n4530) );
  NAND4X1 U9475 ( .A(n4533), .B(n4532), .C(n4531), .D(n4530), .Y(n4537) );
  AOI22X1 U9476 ( .A0(cal_out[436]), .A1(n4910), .B0(cal_out[396]), .B1(n4878), 
        .Y(n4536) );
  AOI222X1 U9477 ( .A0(cal_out[196]), .A1(n4917), .B0(cal_out[276]), .B1(n4881), .C0(cal_out[236]), .C1(n4880), .Y(n4535) );
  AOI22X1 U9478 ( .A0(cal_out[356]), .A1(n4921), .B0(cal_out[156]), .B1(n4883), 
        .Y(n4534) );
  NAND4BXL U9479 ( .AN(n4537), .B(n4536), .C(n4535), .D(n4534), .Y(
        value_out[36]) );
  AOI22X1 U9480 ( .A0(cal_out[515]), .A1(n4894), .B0(cal_out[315]), .B1(n4866), 
        .Y(n4541) );
  AOI22X1 U9481 ( .A0(cal_out[595]), .A1(n4898), .B0(cal_out[555]), .B1(n4868), 
        .Y(n4540) );
  AOI22X1 U9482 ( .A0(cal_out[35]), .A1(n4902), .B0(cal_out[475]), .B1(n4870), 
        .Y(n4539) );
  AOI22X1 U9483 ( .A0(cal_out[115]), .A1(n4906), .B0(cal_out[75]), .B1(n4872), 
        .Y(n4538) );
  NAND4X1 U9484 ( .A(n4541), .B(n4540), .C(n4539), .D(n4538), .Y(n4545) );
  AOI22X1 U9485 ( .A0(cal_out[435]), .A1(n4910), .B0(cal_out[395]), .B1(n4878), 
        .Y(n4544) );
  AOI222X1 U9486 ( .A0(cal_out[195]), .A1(n4917), .B0(cal_out[275]), .B1(n4881), .C0(cal_out[235]), .C1(n4880), .Y(n4543) );
  AOI22X1 U9487 ( .A0(cal_out[355]), .A1(n4921), .B0(cal_out[155]), .B1(n4883), 
        .Y(n4542) );
  NAND4BXL U9488 ( .AN(n4545), .B(n4544), .C(n4543), .D(n4542), .Y(
        value_out[35]) );
  AOI22X1 U9489 ( .A0(cal_out[514]), .A1(n4894), .B0(cal_out[314]), .B1(n4866), 
        .Y(n4549) );
  AOI22X1 U9490 ( .A0(cal_out[594]), .A1(n4898), .B0(cal_out[554]), .B1(n4868), 
        .Y(n4548) );
  AOI22X1 U9491 ( .A0(cal_out[34]), .A1(n4902), .B0(cal_out[474]), .B1(n4870), 
        .Y(n4547) );
  AOI22X1 U9492 ( .A0(cal_out[114]), .A1(n4906), .B0(cal_out[74]), .B1(n4872), 
        .Y(n4546) );
  NAND4X1 U9493 ( .A(n4549), .B(n4548), .C(n4547), .D(n4546), .Y(n4553) );
  AOI22X1 U9494 ( .A0(cal_out[434]), .A1(n4910), .B0(cal_out[394]), .B1(n4878), 
        .Y(n4552) );
  AOI222X1 U9495 ( .A0(cal_out[194]), .A1(n4917), .B0(cal_out[274]), .B1(n4881), .C0(cal_out[234]), .C1(n4880), .Y(n4551) );
  AOI22X1 U9496 ( .A0(cal_out[354]), .A1(n4921), .B0(cal_out[154]), .B1(n4883), 
        .Y(n4550) );
  NAND4BXL U9497 ( .AN(n4553), .B(n4552), .C(n4551), .D(n4550), .Y(
        value_out[34]) );
  AOI22X1 U9498 ( .A0(cal_out[513]), .A1(n4894), .B0(cal_out[313]), .B1(n4866), 
        .Y(n4557) );
  AOI22X1 U9499 ( .A0(cal_out[593]), .A1(n4898), .B0(cal_out[553]), .B1(n4868), 
        .Y(n4556) );
  AOI22X1 U9500 ( .A0(cal_out[33]), .A1(n4902), .B0(cal_out[473]), .B1(n4870), 
        .Y(n4555) );
  AOI22X1 U9501 ( .A0(cal_out[113]), .A1(n4906), .B0(cal_out[73]), .B1(n4872), 
        .Y(n4554) );
  NAND4X1 U9502 ( .A(n4557), .B(n4556), .C(n4555), .D(n4554), .Y(n4561) );
  AOI22X1 U9503 ( .A0(cal_out[433]), .A1(n4910), .B0(cal_out[393]), .B1(n4878), 
        .Y(n4560) );
  AOI222X1 U9504 ( .A0(cal_out[193]), .A1(n4917), .B0(cal_out[273]), .B1(n4881), .C0(cal_out[233]), .C1(n4880), .Y(n4559) );
  AOI22X1 U9505 ( .A0(cal_out[353]), .A1(n4921), .B0(cal_out[153]), .B1(n4883), 
        .Y(n4558) );
  NAND4BXL U9506 ( .AN(n4561), .B(n4560), .C(n4559), .D(n4558), .Y(
        value_out[33]) );
  AOI22X1 U9507 ( .A0(cal_out[512]), .A1(n4894), .B0(cal_out[312]), .B1(n4866), 
        .Y(n4565) );
  AOI22X1 U9508 ( .A0(cal_out[592]), .A1(n4898), .B0(cal_out[552]), .B1(n4868), 
        .Y(n4564) );
  AOI22X1 U9509 ( .A0(cal_out[32]), .A1(n4902), .B0(cal_out[472]), .B1(n4870), 
        .Y(n4563) );
  AOI22X1 U9510 ( .A0(cal_out[112]), .A1(n4906), .B0(cal_out[72]), .B1(n4872), 
        .Y(n4562) );
  NAND4X1 U9511 ( .A(n4565), .B(n4564), .C(n4563), .D(n4562), .Y(n4569) );
  AOI22X1 U9512 ( .A0(cal_out[432]), .A1(n4910), .B0(cal_out[392]), .B1(n4878), 
        .Y(n4568) );
  AOI222X1 U9513 ( .A0(cal_out[192]), .A1(n4917), .B0(cal_out[272]), .B1(n4881), .C0(cal_out[232]), .C1(n4880), .Y(n4567) );
  AOI22X1 U9514 ( .A0(cal_out[352]), .A1(n4921), .B0(cal_out[152]), .B1(n4883), 
        .Y(n4566) );
  NAND4BXL U9515 ( .AN(n4569), .B(n4568), .C(n4567), .D(n4566), .Y(
        value_out[32]) );
  AOI22X1 U9516 ( .A0(cal_out[511]), .A1(n4894), .B0(cal_out[311]), .B1(n4866), 
        .Y(n4573) );
  AOI22X1 U9517 ( .A0(cal_out[591]), .A1(n4898), .B0(cal_out[551]), .B1(n4868), 
        .Y(n4572) );
  AOI22X1 U9518 ( .A0(cal_out[31]), .A1(n4902), .B0(cal_out[471]), .B1(n4870), 
        .Y(n4571) );
  AOI22X1 U9519 ( .A0(cal_out[111]), .A1(n4906), .B0(cal_out[71]), .B1(n4872), 
        .Y(n4570) );
  NAND4X1 U9520 ( .A(n4573), .B(n4572), .C(n4571), .D(n4570), .Y(n4577) );
  AOI22X1 U9521 ( .A0(cal_out[431]), .A1(n4910), .B0(cal_out[391]), .B1(n4878), 
        .Y(n4576) );
  AOI222X1 U9522 ( .A0(cal_out[191]), .A1(n4917), .B0(cal_out[271]), .B1(n4881), .C0(cal_out[231]), .C1(n4880), .Y(n4575) );
  AOI22X1 U9523 ( .A0(cal_out[351]), .A1(n4921), .B0(cal_out[151]), .B1(n4883), 
        .Y(n4574) );
  NAND4BXL U9524 ( .AN(n4577), .B(n4576), .C(n4575), .D(n4574), .Y(
        value_out[31]) );
  AOI22X1 U9525 ( .A0(cal_out[510]), .A1(n4894), .B0(cal_out[310]), .B1(n4866), 
        .Y(n4581) );
  AOI22X1 U9526 ( .A0(cal_out[590]), .A1(n4898), .B0(cal_out[550]), .B1(n4868), 
        .Y(n4580) );
  AOI22X1 U9527 ( .A0(cal_out[30]), .A1(n4902), .B0(cal_out[470]), .B1(n4870), 
        .Y(n4579) );
  AOI22X1 U9528 ( .A0(cal_out[110]), .A1(n4906), .B0(cal_out[70]), .B1(n4872), 
        .Y(n4578) );
  NAND4X1 U9529 ( .A(n4581), .B(n4580), .C(n4579), .D(n4578), .Y(n4585) );
  AOI22X1 U9530 ( .A0(cal_out[430]), .A1(n4910), .B0(cal_out[390]), .B1(n4878), 
        .Y(n4584) );
  AOI222X1 U9531 ( .A0(cal_out[190]), .A1(n4917), .B0(cal_out[270]), .B1(n4881), .C0(cal_out[230]), .C1(n4880), .Y(n4583) );
  AOI22X1 U9532 ( .A0(cal_out[350]), .A1(n4921), .B0(cal_out[150]), .B1(n4883), 
        .Y(n4582) );
  NAND4BXL U9533 ( .AN(n4585), .B(n4584), .C(n4583), .D(n4582), .Y(
        value_out[30]) );
  AOI22X1 U9534 ( .A0(cal_out[509]), .A1(n4894), .B0(cal_out[309]), .B1(n4866), 
        .Y(n4589) );
  AOI22X1 U9535 ( .A0(cal_out[589]), .A1(n4898), .B0(cal_out[549]), .B1(n4868), 
        .Y(n4588) );
  AOI22X1 U9536 ( .A0(cal_out[29]), .A1(n4902), .B0(cal_out[469]), .B1(n4870), 
        .Y(n4587) );
  AOI22X1 U9537 ( .A0(cal_out[109]), .A1(n4906), .B0(cal_out[69]), .B1(n4872), 
        .Y(n4586) );
  NAND4X1 U9538 ( .A(n4589), .B(n4588), .C(n4587), .D(n4586), .Y(n4593) );
  AOI22X1 U9539 ( .A0(cal_out[429]), .A1(n4910), .B0(cal_out[389]), .B1(n4878), 
        .Y(n4592) );
  AOI222X1 U9540 ( .A0(cal_out[189]), .A1(n4917), .B0(cal_out[269]), .B1(n4881), .C0(cal_out[229]), .C1(n4880), .Y(n4591) );
  AOI22X1 U9541 ( .A0(cal_out[349]), .A1(n4921), .B0(cal_out[149]), .B1(n4883), 
        .Y(n4590) );
  NAND4BXL U9542 ( .AN(n4593), .B(n4592), .C(n4591), .D(n4590), .Y(
        value_out[29]) );
  AOI22X1 U9543 ( .A0(cal_out[508]), .A1(n4894), .B0(cal_out[308]), .B1(n4866), 
        .Y(n4597) );
  AOI22X1 U9544 ( .A0(cal_out[588]), .A1(n4898), .B0(cal_out[548]), .B1(n4868), 
        .Y(n4596) );
  AOI22X1 U9545 ( .A0(cal_out[28]), .A1(n4902), .B0(cal_out[468]), .B1(n4870), 
        .Y(n4595) );
  AOI22X1 U9546 ( .A0(cal_out[108]), .A1(n4906), .B0(cal_out[68]), .B1(n4872), 
        .Y(n4594) );
  NAND4X1 U9547 ( .A(n4597), .B(n4596), .C(n4595), .D(n4594), .Y(n4601) );
  AOI22X1 U9548 ( .A0(cal_out[428]), .A1(n4910), .B0(cal_out[388]), .B1(n4878), 
        .Y(n4600) );
  AOI222X1 U9549 ( .A0(cal_out[188]), .A1(n4917), .B0(cal_out[268]), .B1(n4881), .C0(cal_out[228]), .C1(n4880), .Y(n4599) );
  AOI22X1 U9550 ( .A0(cal_out[348]), .A1(n4921), .B0(cal_out[148]), .B1(n4883), 
        .Y(n4598) );
  NAND4BXL U9551 ( .AN(n4601), .B(n4600), .C(n4599), .D(n4598), .Y(
        value_out[28]) );
  AOI22X1 U9552 ( .A0(cal_out[507]), .A1(n4894), .B0(cal_out[307]), .B1(n4866), 
        .Y(n4605) );
  AOI22X1 U9553 ( .A0(cal_out[587]), .A1(n4898), .B0(cal_out[547]), .B1(n4868), 
        .Y(n4604) );
  AOI22X1 U9554 ( .A0(cal_out[27]), .A1(n4902), .B0(cal_out[467]), .B1(n4870), 
        .Y(n4603) );
  AOI22X1 U9555 ( .A0(cal_out[107]), .A1(n4906), .B0(cal_out[67]), .B1(n4872), 
        .Y(n4602) );
  NAND4X1 U9556 ( .A(n4605), .B(n4604), .C(n4603), .D(n4602), .Y(n4609) );
  AOI22X1 U9557 ( .A0(cal_out[427]), .A1(n4910), .B0(cal_out[387]), .B1(n4878), 
        .Y(n4608) );
  AOI222X1 U9558 ( .A0(cal_out[187]), .A1(n4917), .B0(cal_out[267]), .B1(n4881), .C0(cal_out[227]), .C1(n4880), .Y(n4607) );
  AOI22X1 U9559 ( .A0(cal_out[347]), .A1(n4921), .B0(cal_out[147]), .B1(n4883), 
        .Y(n4606) );
  NAND4BXL U9560 ( .AN(n4609), .B(n4608), .C(n4607), .D(n4606), .Y(
        value_out[27]) );
  AOI22X1 U9561 ( .A0(cal_out[506]), .A1(n4867), .B0(cal_out[306]), .B1(n4866), 
        .Y(n4613) );
  AOI22X1 U9562 ( .A0(cal_out[586]), .A1(n4869), .B0(cal_out[546]), .B1(n4868), 
        .Y(n4612) );
  AOI22X1 U9563 ( .A0(cal_out[26]), .A1(n4871), .B0(cal_out[466]), .B1(n4870), 
        .Y(n4611) );
  AOI22X1 U9564 ( .A0(cal_out[106]), .A1(n4873), .B0(cal_out[66]), .B1(n4872), 
        .Y(n4610) );
  NAND4X1 U9565 ( .A(n4613), .B(n4612), .C(n4611), .D(n4610), .Y(n4617) );
  AOI22X1 U9566 ( .A0(cal_out[426]), .A1(n4879), .B0(cal_out[386]), .B1(n4878), 
        .Y(n4616) );
  AOI222X1 U9567 ( .A0(cal_out[186]), .A1(n4882), .B0(cal_out[266]), .B1(n4881), .C0(cal_out[226]), .C1(n4880), .Y(n4615) );
  AOI22X1 U9568 ( .A0(cal_out[346]), .A1(n4884), .B0(cal_out[146]), .B1(n4883), 
        .Y(n4614) );
  NAND4BXL U9569 ( .AN(n4617), .B(n4616), .C(n4615), .D(n4614), .Y(
        value_out[26]) );
  AOI22X1 U9570 ( .A0(cal_out[505]), .A1(n4867), .B0(cal_out[305]), .B1(n4866), 
        .Y(n4621) );
  AOI22X1 U9571 ( .A0(cal_out[585]), .A1(n4869), .B0(cal_out[545]), .B1(n4868), 
        .Y(n4620) );
  AOI22X1 U9572 ( .A0(cal_out[25]), .A1(n4871), .B0(cal_out[465]), .B1(n4870), 
        .Y(n4619) );
  AOI22X1 U9573 ( .A0(cal_out[105]), .A1(n4873), .B0(cal_out[65]), .B1(n4872), 
        .Y(n4618) );
  NAND4X1 U9574 ( .A(n4621), .B(n4620), .C(n4619), .D(n4618), .Y(n4625) );
  AOI22X1 U9575 ( .A0(cal_out[425]), .A1(n4879), .B0(cal_out[385]), .B1(n4878), 
        .Y(n4624) );
  AOI222X1 U9576 ( .A0(cal_out[185]), .A1(n4882), .B0(cal_out[265]), .B1(n4914), .C0(cal_out[225]), .C1(n4880), .Y(n4623) );
  AOI22X1 U9577 ( .A0(cal_out[345]), .A1(n4884), .B0(cal_out[145]), .B1(n4883), 
        .Y(n4622) );
  NAND4BXL U9578 ( .AN(n4625), .B(n4624), .C(n4623), .D(n4622), .Y(
        value_out[25]) );
  AOI22X1 U9579 ( .A0(cal_out[504]), .A1(n4867), .B0(cal_out[304]), .B1(n4866), 
        .Y(n4629) );
  AOI22X1 U9580 ( .A0(cal_out[584]), .A1(n4869), .B0(cal_out[544]), .B1(n4868), 
        .Y(n4628) );
  AOI22X1 U9581 ( .A0(cal_out[24]), .A1(n4871), .B0(cal_out[464]), .B1(n4870), 
        .Y(n4627) );
  AOI22X1 U9582 ( .A0(cal_out[104]), .A1(n4873), .B0(cal_out[64]), .B1(n4872), 
        .Y(n4626) );
  NAND4X1 U9583 ( .A(n4629), .B(n4628), .C(n4627), .D(n4626), .Y(n4633) );
  AOI22X1 U9584 ( .A0(cal_out[424]), .A1(n4879), .B0(cal_out[384]), .B1(n4878), 
        .Y(n4632) );
  AOI222X1 U9585 ( .A0(cal_out[184]), .A1(n4882), .B0(cal_out[264]), .B1(n4881), .C0(cal_out[224]), .C1(n4880), .Y(n4631) );
  AOI22X1 U9586 ( .A0(cal_out[344]), .A1(n4884), .B0(cal_out[144]), .B1(n4883), 
        .Y(n4630) );
  NAND4BXL U9587 ( .AN(n4633), .B(n4632), .C(n4631), .D(n4630), .Y(
        value_out[24]) );
  AOI22X1 U9588 ( .A0(cal_out[503]), .A1(n4867), .B0(cal_out[303]), .B1(n4866), 
        .Y(n4637) );
  AOI22X1 U9589 ( .A0(cal_out[583]), .A1(n4869), .B0(cal_out[543]), .B1(n4868), 
        .Y(n4636) );
  AOI22X1 U9590 ( .A0(cal_out[23]), .A1(n4871), .B0(cal_out[463]), .B1(n4870), 
        .Y(n4635) );
  AOI22X1 U9591 ( .A0(cal_out[103]), .A1(n4873), .B0(cal_out[63]), .B1(n4872), 
        .Y(n4634) );
  NAND4X1 U9592 ( .A(n4637), .B(n4636), .C(n4635), .D(n4634), .Y(n4641) );
  AOI22X1 U9593 ( .A0(cal_out[423]), .A1(n4879), .B0(cal_out[383]), .B1(n4878), 
        .Y(n4640) );
  AOI222X1 U9594 ( .A0(cal_out[183]), .A1(n4882), .B0(cal_out[263]), .B1(n4881), .C0(cal_out[223]), .C1(n4880), .Y(n4639) );
  AOI22X1 U9595 ( .A0(cal_out[343]), .A1(n4884), .B0(cal_out[143]), .B1(n4883), 
        .Y(n4638) );
  NAND4BXL U9596 ( .AN(n4641), .B(n4640), .C(n4639), .D(n4638), .Y(
        value_out[23]) );
  AOI22X1 U9597 ( .A0(cal_out[502]), .A1(n4867), .B0(cal_out[302]), .B1(n4866), 
        .Y(n4645) );
  AOI22X1 U9598 ( .A0(cal_out[582]), .A1(n4869), .B0(cal_out[542]), .B1(n4868), 
        .Y(n4644) );
  AOI22X1 U9599 ( .A0(cal_out[22]), .A1(n4871), .B0(cal_out[462]), .B1(n4870), 
        .Y(n4643) );
  AOI22X1 U9600 ( .A0(cal_out[102]), .A1(n4873), .B0(cal_out[62]), .B1(n4872), 
        .Y(n4642) );
  NAND4X1 U9601 ( .A(n4645), .B(n4644), .C(n4643), .D(n4642), .Y(n4649) );
  AOI22X1 U9602 ( .A0(cal_out[422]), .A1(n4879), .B0(cal_out[382]), .B1(n4878), 
        .Y(n4648) );
  AOI222X1 U9603 ( .A0(cal_out[182]), .A1(n4882), .B0(cal_out[262]), .B1(n4881), .C0(cal_out[222]), .C1(n4880), .Y(n4647) );
  AOI22X1 U9604 ( .A0(cal_out[342]), .A1(n4884), .B0(cal_out[142]), .B1(n4883), 
        .Y(n4646) );
  NAND4BXL U9605 ( .AN(n4649), .B(n4648), .C(n4647), .D(n4646), .Y(
        value_out[22]) );
  AOI22X1 U9606 ( .A0(cal_out[501]), .A1(n4867), .B0(cal_out[301]), .B1(n4866), 
        .Y(n4653) );
  AOI22X1 U9607 ( .A0(cal_out[581]), .A1(n4869), .B0(cal_out[541]), .B1(n4868), 
        .Y(n4652) );
  AOI22X1 U9608 ( .A0(cal_out[21]), .A1(n4871), .B0(cal_out[461]), .B1(n4870), 
        .Y(n4651) );
  AOI22X1 U9609 ( .A0(cal_out[101]), .A1(n4873), .B0(cal_out[61]), .B1(n4872), 
        .Y(n4650) );
  NAND4X1 U9610 ( .A(n4653), .B(n4652), .C(n4651), .D(n4650), .Y(n4657) );
  AOI22X1 U9611 ( .A0(cal_out[421]), .A1(n4879), .B0(cal_out[381]), .B1(n4878), 
        .Y(n4656) );
  AOI222X1 U9612 ( .A0(cal_out[181]), .A1(n4882), .B0(cal_out[261]), .B1(n4914), .C0(cal_out[221]), .C1(n4880), .Y(n4655) );
  AOI22X1 U9613 ( .A0(cal_out[341]), .A1(n4884), .B0(cal_out[141]), .B1(n4883), 
        .Y(n4654) );
  NAND4BXL U9614 ( .AN(n4657), .B(n4656), .C(n4655), .D(n4654), .Y(
        value_out[21]) );
  AOI22X1 U9615 ( .A0(cal_out[500]), .A1(n4867), .B0(cal_out[300]), .B1(n4866), 
        .Y(n4661) );
  AOI22X1 U9616 ( .A0(cal_out[580]), .A1(n4869), .B0(cal_out[540]), .B1(n4868), 
        .Y(n4660) );
  AOI22X1 U9617 ( .A0(cal_out[20]), .A1(n4871), .B0(cal_out[460]), .B1(n4870), 
        .Y(n4659) );
  AOI22X1 U9618 ( .A0(cal_out[100]), .A1(n4873), .B0(cal_out[60]), .B1(n4872), 
        .Y(n4658) );
  NAND4X1 U9619 ( .A(n4661), .B(n4660), .C(n4659), .D(n4658), .Y(n4665) );
  AOI22X1 U9620 ( .A0(cal_out[420]), .A1(n4879), .B0(cal_out[380]), .B1(n4878), 
        .Y(n4664) );
  AOI222X1 U9621 ( .A0(cal_out[180]), .A1(n4882), .B0(cal_out[260]), .B1(n4881), .C0(cal_out[220]), .C1(n4880), .Y(n4663) );
  AOI22X1 U9622 ( .A0(cal_out[340]), .A1(n4884), .B0(cal_out[140]), .B1(n4883), 
        .Y(n4662) );
  NAND4BXL U9623 ( .AN(n4665), .B(n4664), .C(n4663), .D(n4662), .Y(
        value_out[20]) );
  AOI22X1 U9624 ( .A0(cal_out[499]), .A1(n4867), .B0(cal_out[299]), .B1(n4866), 
        .Y(n4669) );
  AOI22X1 U9625 ( .A0(cal_out[579]), .A1(n4869), .B0(cal_out[539]), .B1(n4868), 
        .Y(n4668) );
  AOI22X1 U9626 ( .A0(cal_out[19]), .A1(n4871), .B0(cal_out[459]), .B1(n4870), 
        .Y(n4667) );
  AOI22X1 U9627 ( .A0(cal_out[99]), .A1(n4873), .B0(cal_out[59]), .B1(n4872), 
        .Y(n4666) );
  NAND4X1 U9628 ( .A(n4669), .B(n4668), .C(n4667), .D(n4666), .Y(n4673) );
  AOI22X1 U9629 ( .A0(cal_out[419]), .A1(n4879), .B0(cal_out[379]), .B1(n4878), 
        .Y(n4672) );
  AOI222X1 U9630 ( .A0(cal_out[179]), .A1(n4882), .B0(cal_out[259]), .B1(n4914), .C0(cal_out[219]), .C1(n4880), .Y(n4671) );
  AOI22X1 U9631 ( .A0(cal_out[339]), .A1(n4884), .B0(cal_out[139]), .B1(n4883), 
        .Y(n4670) );
  NAND4BXL U9632 ( .AN(n4673), .B(n4672), .C(n4671), .D(n4670), .Y(
        value_out[19]) );
  AOI22X1 U9633 ( .A0(cal_out[498]), .A1(n4894), .B0(cal_out[298]), .B1(n4866), 
        .Y(n4677) );
  AOI22X1 U9634 ( .A0(cal_out[578]), .A1(n4898), .B0(cal_out[538]), .B1(n4868), 
        .Y(n4676) );
  AOI22X1 U9635 ( .A0(cal_out[18]), .A1(n4871), .B0(cal_out[458]), .B1(n4870), 
        .Y(n4675) );
  AOI22X1 U9636 ( .A0(cal_out[98]), .A1(n4906), .B0(cal_out[58]), .B1(n4872), 
        .Y(n4674) );
  NAND4X1 U9637 ( .A(n4677), .B(n4676), .C(n4675), .D(n4674), .Y(n4681) );
  AOI22X1 U9638 ( .A0(cal_out[418]), .A1(n4910), .B0(cal_out[378]), .B1(n4878), 
        .Y(n4680) );
  AOI222X1 U9639 ( .A0(cal_out[178]), .A1(n4882), .B0(cal_out[258]), .B1(n4914), .C0(cal_out[218]), .C1(n4880), .Y(n4679) );
  AOI22X1 U9640 ( .A0(cal_out[338]), .A1(n4921), .B0(cal_out[138]), .B1(n4883), 
        .Y(n4678) );
  NAND4BXL U9641 ( .AN(n4681), .B(n4680), .C(n4679), .D(n4678), .Y(
        value_out[18]) );
  AOI22X1 U9642 ( .A0(cal_out[497]), .A1(n4867), .B0(cal_out[297]), .B1(n4866), 
        .Y(n4685) );
  AOI22X1 U9643 ( .A0(cal_out[577]), .A1(n4869), .B0(cal_out[537]), .B1(n4868), 
        .Y(n4684) );
  AOI22X1 U9644 ( .A0(cal_out[17]), .A1(n4871), .B0(cal_out[457]), .B1(n4870), 
        .Y(n4683) );
  AOI22X1 U9645 ( .A0(cal_out[97]), .A1(n4873), .B0(cal_out[57]), .B1(n4872), 
        .Y(n4682) );
  NAND4X1 U9646 ( .A(n4685), .B(n4684), .C(n4683), .D(n4682), .Y(n4689) );
  AOI22X1 U9647 ( .A0(cal_out[417]), .A1(n4879), .B0(cal_out[377]), .B1(n4878), 
        .Y(n4688) );
  AOI222X1 U9648 ( .A0(cal_out[177]), .A1(n4882), .B0(cal_out[257]), .B1(n4881), .C0(cal_out[217]), .C1(n4880), .Y(n4687) );
  AOI22X1 U9649 ( .A0(cal_out[337]), .A1(n4884), .B0(cal_out[137]), .B1(n4883), 
        .Y(n4686) );
  NAND4BXL U9650 ( .AN(n4689), .B(n4688), .C(n4687), .D(n4686), .Y(
        value_out[17]) );
  AOI22X1 U9651 ( .A0(cal_out[496]), .A1(n4867), .B0(cal_out[296]), .B1(n4866), 
        .Y(n4693) );
  AOI22X1 U9652 ( .A0(cal_out[576]), .A1(n4869), .B0(cal_out[536]), .B1(n4868), 
        .Y(n4692) );
  AOI22X1 U9653 ( .A0(cal_out[16]), .A1(n4871), .B0(cal_out[456]), .B1(n4870), 
        .Y(n4691) );
  AOI22X1 U9654 ( .A0(cal_out[96]), .A1(n4873), .B0(cal_out[56]), .B1(n4872), 
        .Y(n4690) );
  NAND4X1 U9655 ( .A(n4693), .B(n4692), .C(n4691), .D(n4690), .Y(n4697) );
  AOI22X1 U9656 ( .A0(cal_out[416]), .A1(n4879), .B0(cal_out[376]), .B1(n4878), 
        .Y(n4696) );
  AOI222X1 U9657 ( .A0(cal_out[176]), .A1(n4882), .B0(cal_out[256]), .B1(n4881), .C0(cal_out[216]), .C1(n4880), .Y(n4695) );
  AOI22X1 U9658 ( .A0(cal_out[336]), .A1(n4884), .B0(cal_out[136]), .B1(n4883), 
        .Y(n4694) );
  NAND4BXL U9659 ( .AN(n4697), .B(n4696), .C(n4695), .D(n4694), .Y(
        value_out[16]) );
  AOI22X1 U9660 ( .A0(cal_out[495]), .A1(n4867), .B0(cal_out[295]), .B1(n4866), 
        .Y(n4701) );
  AOI22X1 U9661 ( .A0(cal_out[575]), .A1(n4869), .B0(cal_out[535]), .B1(n4868), 
        .Y(n4700) );
  AOI22X1 U9662 ( .A0(cal_out[15]), .A1(n4871), .B0(cal_out[455]), .B1(n4870), 
        .Y(n4699) );
  AOI22X1 U9663 ( .A0(cal_out[95]), .A1(n4873), .B0(cal_out[55]), .B1(n4872), 
        .Y(n4698) );
  NAND4X1 U9664 ( .A(n4701), .B(n4700), .C(n4699), .D(n4698), .Y(n4705) );
  AOI22X1 U9665 ( .A0(cal_out[415]), .A1(n4879), .B0(cal_out[375]), .B1(n4878), 
        .Y(n4704) );
  AOI222X1 U9666 ( .A0(cal_out[175]), .A1(n4882), .B0(cal_out[255]), .B1(n4914), .C0(cal_out[215]), .C1(n4912), .Y(n4703) );
  AOI22X1 U9667 ( .A0(cal_out[335]), .A1(n4884), .B0(cal_out[135]), .B1(n4883), 
        .Y(n4702) );
  NAND4BXL U9668 ( .AN(n4705), .B(n4704), .C(n4703), .D(n4702), .Y(
        value_out[15]) );
  AOI22X1 U9669 ( .A0(cal_out[494]), .A1(n4867), .B0(cal_out[294]), .B1(n4866), 
        .Y(n4709) );
  AOI22X1 U9670 ( .A0(cal_out[574]), .A1(n4869), .B0(cal_out[534]), .B1(n4868), 
        .Y(n4708) );
  AOI22X1 U9671 ( .A0(cal_out[14]), .A1(n4871), .B0(cal_out[454]), .B1(n4870), 
        .Y(n4707) );
  AOI22X1 U9672 ( .A0(cal_out[94]), .A1(n4873), .B0(cal_out[54]), .B1(n4872), 
        .Y(n4706) );
  NAND4X1 U9673 ( .A(n4709), .B(n4708), .C(n4707), .D(n4706), .Y(n4713) );
  AOI22X1 U9674 ( .A0(cal_out[414]), .A1(n4879), .B0(cal_out[374]), .B1(n4878), 
        .Y(n4712) );
  AOI222X1 U9675 ( .A0(cal_out[174]), .A1(n4882), .B0(cal_out[254]), .B1(n4914), .C0(cal_out[214]), .C1(n4912), .Y(n4711) );
  AOI22X1 U9676 ( .A0(cal_out[334]), .A1(n4884), .B0(cal_out[134]), .B1(n4883), 
        .Y(n4710) );
  NAND4BXL U9677 ( .AN(n4713), .B(n4712), .C(n4711), .D(n4710), .Y(
        value_out[14]) );
  AOI22X1 U9678 ( .A0(cal_out[493]), .A1(n4867), .B0(cal_out[293]), .B1(n4892), 
        .Y(n4717) );
  AOI22X1 U9679 ( .A0(cal_out[573]), .A1(n4869), .B0(cal_out[533]), .B1(n4896), 
        .Y(n4716) );
  AOI22X1 U9680 ( .A0(cal_out[13]), .A1(n4871), .B0(cal_out[453]), .B1(n4900), 
        .Y(n4715) );
  AOI22X1 U9681 ( .A0(cal_out[93]), .A1(n4873), .B0(cal_out[53]), .B1(n4904), 
        .Y(n4714) );
  NAND4X1 U9682 ( .A(n4717), .B(n4716), .C(n4715), .D(n4714), .Y(n4721) );
  AOI22X1 U9683 ( .A0(cal_out[413]), .A1(n4879), .B0(cal_out[373]), .B1(n4908), 
        .Y(n4720) );
  AOI222X1 U9684 ( .A0(cal_out[173]), .A1(n4916), .B0(cal_out[253]), .B1(n4914), .C0(cal_out[213]), .C1(n4880), .Y(n4719) );
  AOI22X1 U9685 ( .A0(cal_out[333]), .A1(n4884), .B0(cal_out[133]), .B1(n4919), 
        .Y(n4718) );
  NAND4BXL U9686 ( .AN(n4721), .B(n4720), .C(n4719), .D(n4718), .Y(
        value_out[13]) );
  AOI22X1 U9687 ( .A0(cal_out[492]), .A1(n4894), .B0(cal_out[292]), .B1(n4892), 
        .Y(n4725) );
  AOI22X1 U9688 ( .A0(cal_out[572]), .A1(n4898), .B0(cal_out[532]), .B1(n4896), 
        .Y(n4724) );
  AOI22X1 U9689 ( .A0(cal_out[12]), .A1(n4902), .B0(cal_out[452]), .B1(n4900), 
        .Y(n4723) );
  AOI22X1 U9690 ( .A0(cal_out[92]), .A1(n4906), .B0(cal_out[52]), .B1(n4904), 
        .Y(n4722) );
  NAND4X1 U9691 ( .A(n4725), .B(n4724), .C(n4723), .D(n4722), .Y(n4729) );
  AOI22X1 U9692 ( .A0(cal_out[412]), .A1(n4910), .B0(cal_out[372]), .B1(n4908), 
        .Y(n4728) );
  AOI222X1 U9693 ( .A0(cal_out[172]), .A1(n4916), .B0(cal_out[252]), .B1(n4914), .C0(cal_out[212]), .C1(n4880), .Y(n4727) );
  AOI22X1 U9694 ( .A0(cal_out[332]), .A1(n4921), .B0(cal_out[132]), .B1(n4919), 
        .Y(n4726) );
  NAND4BXL U9695 ( .AN(n4729), .B(n4728), .C(n4727), .D(n4726), .Y(
        value_out[12]) );
  AOI22X1 U9696 ( .A0(cal_out[491]), .A1(n4867), .B0(cal_out[291]), .B1(n4892), 
        .Y(n4733) );
  AOI22X1 U9697 ( .A0(cal_out[571]), .A1(n4869), .B0(cal_out[531]), .B1(n4896), 
        .Y(n4732) );
  AOI22X1 U9698 ( .A0(cal_out[11]), .A1(n4871), .B0(cal_out[451]), .B1(n4900), 
        .Y(n4731) );
  AOI22X1 U9699 ( .A0(cal_out[91]), .A1(n4873), .B0(cal_out[51]), .B1(n4904), 
        .Y(n4730) );
  NAND4X1 U9700 ( .A(n4733), .B(n4732), .C(n4731), .D(n4730), .Y(n4737) );
  AOI22X1 U9701 ( .A0(cal_out[411]), .A1(n4879), .B0(cal_out[371]), .B1(n4908), 
        .Y(n4736) );
  AOI222X1 U9702 ( .A0(cal_out[171]), .A1(n4916), .B0(cal_out[251]), .B1(n4914), .C0(cal_out[211]), .C1(n4880), .Y(n4735) );
  AOI22X1 U9703 ( .A0(cal_out[331]), .A1(n4884), .B0(cal_out[131]), .B1(n4919), 
        .Y(n4734) );
  NAND4BXL U9704 ( .AN(n4737), .B(n4736), .C(n4735), .D(n4734), .Y(
        value_out[11]) );
  AOI22X1 U9705 ( .A0(cal_out[490]), .A1(n4867), .B0(cal_out[290]), .B1(n4892), 
        .Y(n4741) );
  AOI22X1 U9706 ( .A0(cal_out[570]), .A1(n4869), .B0(cal_out[530]), .B1(n4896), 
        .Y(n4740) );
  AOI22X1 U9707 ( .A0(cal_out[10]), .A1(n4871), .B0(cal_out[450]), .B1(n4900), 
        .Y(n4739) );
  AOI22X1 U9708 ( .A0(cal_out[90]), .A1(n4873), .B0(cal_out[50]), .B1(n4904), 
        .Y(n4738) );
  NAND4X1 U9709 ( .A(n4741), .B(n4740), .C(n4739), .D(n4738), .Y(n4745) );
  AOI22X1 U9710 ( .A0(cal_out[410]), .A1(n4879), .B0(cal_out[370]), .B1(n4908), 
        .Y(n4744) );
  AOI222X1 U9711 ( .A0(cal_out[170]), .A1(n4916), .B0(cal_out[250]), .B1(n4914), .C0(cal_out[210]), .C1(n4880), .Y(n4743) );
  AOI22X1 U9712 ( .A0(cal_out[330]), .A1(n4884), .B0(cal_out[130]), .B1(n4919), 
        .Y(n4742) );
  NAND4BXL U9713 ( .AN(n4745), .B(n4744), .C(n4743), .D(n4742), .Y(
        value_out[10]) );
  AOI22X1 U9714 ( .A0(cal_out[489]), .A1(n4867), .B0(cal_out[289]), .B1(n4892), 
        .Y(n4749) );
  AOI22X1 U9715 ( .A0(cal_out[569]), .A1(n4869), .B0(cal_out[529]), .B1(n4896), 
        .Y(n4748) );
  AOI22X1 U9716 ( .A0(cal_out[9]), .A1(n4871), .B0(cal_out[449]), .B1(n4900), 
        .Y(n4747) );
  AOI22X1 U9717 ( .A0(cal_out[89]), .A1(n4873), .B0(cal_out[49]), .B1(n4904), 
        .Y(n4746) );
  NAND4X1 U9718 ( .A(n4749), .B(n4748), .C(n4747), .D(n4746), .Y(n4753) );
  AOI22X1 U9719 ( .A0(cal_out[409]), .A1(n4879), .B0(cal_out[369]), .B1(n4908), 
        .Y(n4752) );
  AOI222X1 U9720 ( .A0(cal_out[169]), .A1(n4916), .B0(cal_out[249]), .B1(n4914), .C0(cal_out[209]), .C1(n4912), .Y(n4751) );
  AOI22X1 U9721 ( .A0(cal_out[329]), .A1(n4884), .B0(cal_out[129]), .B1(n4919), 
        .Y(n4750) );
  NAND4BXL U9722 ( .AN(n4753), .B(n4752), .C(n4751), .D(n4750), .Y(
        value_out[9]) );
  AOI22X1 U9723 ( .A0(cal_out[488]), .A1(n4894), .B0(cal_out[288]), .B1(n4892), 
        .Y(n4757) );
  AOI22X1 U9724 ( .A0(cal_out[568]), .A1(n4898), .B0(cal_out[528]), .B1(n4896), 
        .Y(n4756) );
  AOI22X1 U9725 ( .A0(cal_out[8]), .A1(n4902), .B0(cal_out[448]), .B1(n4900), 
        .Y(n4755) );
  AOI22X1 U9726 ( .A0(cal_out[88]), .A1(n4906), .B0(cal_out[48]), .B1(n4904), 
        .Y(n4754) );
  NAND4X1 U9727 ( .A(n4757), .B(n4756), .C(n4755), .D(n4754), .Y(n4761) );
  AOI22X1 U9728 ( .A0(cal_out[408]), .A1(n4910), .B0(cal_out[368]), .B1(n4908), 
        .Y(n4760) );
  AOI222X1 U9729 ( .A0(cal_out[168]), .A1(n4916), .B0(cal_out[248]), .B1(n4914), .C0(cal_out[208]), .C1(n4880), .Y(n4759) );
  AOI22X1 U9730 ( .A0(cal_out[328]), .A1(n4921), .B0(cal_out[128]), .B1(n4919), 
        .Y(n4758) );
  NAND4BXL U9731 ( .AN(n4761), .B(n4760), .C(n4759), .D(n4758), .Y(
        value_out[8]) );
  AOI22X1 U9732 ( .A0(cal_out[487]), .A1(n4867), .B0(cal_out[287]), .B1(n4892), 
        .Y(n4765) );
  AOI22X1 U9733 ( .A0(cal_out[567]), .A1(n4869), .B0(cal_out[527]), .B1(n4896), 
        .Y(n4764) );
  AOI22X1 U9734 ( .A0(cal_out[7]), .A1(n4871), .B0(cal_out[447]), .B1(n4900), 
        .Y(n4763) );
  AOI22X1 U9735 ( .A0(cal_out[87]), .A1(n4873), .B0(cal_out[47]), .B1(n4904), 
        .Y(n4762) );
  NAND4X1 U9736 ( .A(n4765), .B(n4764), .C(n4763), .D(n4762), .Y(n4769) );
  AOI22X1 U9737 ( .A0(cal_out[407]), .A1(n4879), .B0(cal_out[367]), .B1(n4908), 
        .Y(n4768) );
  AOI222X1 U9738 ( .A0(cal_out[167]), .A1(n4916), .B0(cal_out[247]), .B1(n4914), .C0(cal_out[207]), .C1(n4912), .Y(n4767) );
  AOI22X1 U9739 ( .A0(cal_out[327]), .A1(n4884), .B0(cal_out[127]), .B1(n4919), 
        .Y(n4766) );
  NAND4BXL U9740 ( .AN(n4769), .B(n4768), .C(n4767), .D(n4766), .Y(
        value_out[7]) );
  AOI22X1 U9741 ( .A0(cal_out[486]), .A1(n4867), .B0(cal_out[286]), .B1(n4892), 
        .Y(n4773) );
  AOI22X1 U9742 ( .A0(cal_out[566]), .A1(n4869), .B0(cal_out[526]), .B1(n4896), 
        .Y(n4772) );
  AOI22X1 U9743 ( .A0(cal_out[6]), .A1(n4871), .B0(cal_out[446]), .B1(n4900), 
        .Y(n4771) );
  AOI22X1 U9744 ( .A0(cal_out[86]), .A1(n4873), .B0(cal_out[46]), .B1(n4904), 
        .Y(n4770) );
  NAND4X1 U9745 ( .A(n4773), .B(n4772), .C(n4771), .D(n4770), .Y(n4777) );
  AOI22X1 U9746 ( .A0(cal_out[406]), .A1(n4879), .B0(cal_out[366]), .B1(n4908), 
        .Y(n4776) );
  AOI222X1 U9747 ( .A0(cal_out[166]), .A1(n4916), .B0(cal_out[246]), .B1(n4914), .C0(cal_out[206]), .C1(n4912), .Y(n4775) );
  AOI22X1 U9748 ( .A0(cal_out[326]), .A1(n4884), .B0(cal_out[126]), .B1(n4919), 
        .Y(n4774) );
  NAND4BXL U9749 ( .AN(n4777), .B(n4776), .C(n4775), .D(n4774), .Y(
        value_out[6]) );
  AOI22X1 U9750 ( .A0(cal_out[485]), .A1(n4867), .B0(cal_out[285]), .B1(n4892), 
        .Y(n4781) );
  AOI22X1 U9751 ( .A0(cal_out[565]), .A1(n4869), .B0(cal_out[525]), .B1(n4896), 
        .Y(n4780) );
  AOI22X1 U9752 ( .A0(cal_out[5]), .A1(n4871), .B0(cal_out[445]), .B1(n4900), 
        .Y(n4779) );
  AOI22X1 U9753 ( .A0(cal_out[85]), .A1(n4873), .B0(cal_out[45]), .B1(n4904), 
        .Y(n4778) );
  NAND4X1 U9754 ( .A(n4781), .B(n4780), .C(n4779), .D(n4778), .Y(n4785) );
  AOI22X1 U9755 ( .A0(cal_out[405]), .A1(n4879), .B0(cal_out[365]), .B1(n4908), 
        .Y(n4784) );
  AOI222X1 U9756 ( .A0(cal_out[165]), .A1(n4916), .B0(cal_out[245]), .B1(n4914), .C0(cal_out[205]), .C1(n4880), .Y(n4783) );
  AOI22X1 U9757 ( .A0(cal_out[325]), .A1(n4884), .B0(cal_out[125]), .B1(n4919), 
        .Y(n4782) );
  NAND4BXL U9758 ( .AN(n4785), .B(n4784), .C(n4783), .D(n4782), .Y(
        value_out[5]) );
  AOI22X1 U9759 ( .A0(cal_out[484]), .A1(n4894), .B0(cal_out[284]), .B1(n4892), 
        .Y(n4789) );
  AOI22X1 U9760 ( .A0(cal_out[564]), .A1(n4898), .B0(cal_out[524]), .B1(n4896), 
        .Y(n4788) );
  AOI22X1 U9761 ( .A0(cal_out[4]), .A1(n4902), .B0(cal_out[444]), .B1(n4900), 
        .Y(n4787) );
  AOI22X1 U9762 ( .A0(cal_out[84]), .A1(n4906), .B0(cal_out[44]), .B1(n4904), 
        .Y(n4786) );
  NAND4X1 U9763 ( .A(n4789), .B(n4788), .C(n4787), .D(n4786), .Y(n4793) );
  AOI22X1 U9764 ( .A0(cal_out[404]), .A1(n4910), .B0(cal_out[364]), .B1(n4908), 
        .Y(n4792) );
  AOI222X1 U9765 ( .A0(cal_out[164]), .A1(n4916), .B0(cal_out[244]), .B1(n4914), .C0(cal_out[204]), .C1(n4912), .Y(n4791) );
  AOI22X1 U9766 ( .A0(cal_out[324]), .A1(n4921), .B0(cal_out[124]), .B1(n4919), 
        .Y(n4790) );
  NAND4BXL U9767 ( .AN(n4793), .B(n4792), .C(n4791), .D(n4790), .Y(
        value_out[4]) );
  AOI22X1 U9768 ( .A0(cal_out[483]), .A1(n4867), .B0(cal_out[283]), .B1(n4892), 
        .Y(n4797) );
  AOI22X1 U9769 ( .A0(cal_out[563]), .A1(n4869), .B0(cal_out[523]), .B1(n4896), 
        .Y(n4796) );
  AOI22X1 U9770 ( .A0(cal_out[3]), .A1(n4871), .B0(cal_out[443]), .B1(n4900), 
        .Y(n4795) );
  AOI22X1 U9771 ( .A0(cal_out[83]), .A1(n4873), .B0(cal_out[43]), .B1(n4904), 
        .Y(n4794) );
  NAND4X1 U9772 ( .A(n4797), .B(n4796), .C(n4795), .D(n4794), .Y(n4801) );
  AOI22X1 U9773 ( .A0(cal_out[403]), .A1(n4879), .B0(cal_out[363]), .B1(n4908), 
        .Y(n4800) );
  AOI222X1 U9774 ( .A0(cal_out[163]), .A1(n4916), .B0(cal_out[243]), .B1(n4881), .C0(cal_out[203]), .C1(n4912), .Y(n4799) );
  AOI22X1 U9775 ( .A0(cal_out[323]), .A1(n4884), .B0(cal_out[123]), .B1(n4919), 
        .Y(n4798) );
  NAND4BXL U9776 ( .AN(n4801), .B(n4800), .C(n4799), .D(n4798), .Y(
        value_out[3]) );
  AOI22X1 U9777 ( .A0(cal_out[482]), .A1(n4867), .B0(cal_out[282]), .B1(n4892), 
        .Y(n4805) );
  AOI22X1 U9778 ( .A0(cal_out[562]), .A1(n4869), .B0(cal_out[522]), .B1(n4896), 
        .Y(n4804) );
  AOI22X1 U9779 ( .A0(cal_out[2]), .A1(n4871), .B0(cal_out[442]), .B1(n4900), 
        .Y(n4803) );
  AOI22X1 U9780 ( .A0(cal_out[82]), .A1(n4873), .B0(cal_out[42]), .B1(n4904), 
        .Y(n4802) );
  NAND4X1 U9781 ( .A(n4805), .B(n4804), .C(n4803), .D(n4802), .Y(n4809) );
  AOI22X1 U9782 ( .A0(cal_out[402]), .A1(n4879), .B0(cal_out[362]), .B1(n4908), 
        .Y(n4808) );
  AOI222X1 U9783 ( .A0(cal_out[162]), .A1(n4916), .B0(cal_out[242]), .B1(n4881), .C0(cal_out[202]), .C1(n4912), .Y(n4807) );
  AOI22X1 U9784 ( .A0(cal_out[322]), .A1(n4884), .B0(cal_out[122]), .B1(n4919), 
        .Y(n4806) );
  NAND4BXL U9785 ( .AN(n4809), .B(n4808), .C(n4807), .D(n4806), .Y(
        value_out[2]) );
  AOI22X1 U9786 ( .A0(cal_out[481]), .A1(n4867), .B0(cal_out[281]), .B1(n4892), 
        .Y(n4813) );
  AOI22X1 U9787 ( .A0(cal_out[561]), .A1(n4869), .B0(cal_out[521]), .B1(n4896), 
        .Y(n4812) );
  AOI22X1 U9788 ( .A0(cal_out[1]), .A1(n4871), .B0(cal_out[441]), .B1(n4900), 
        .Y(n4811) );
  AOI22X1 U9789 ( .A0(cal_out[81]), .A1(n4873), .B0(cal_out[41]), .B1(n4904), 
        .Y(n4810) );
  NAND4X1 U9790 ( .A(n4813), .B(n4812), .C(n4811), .D(n4810), .Y(n4817) );
  AOI22X1 U9791 ( .A0(cal_out[401]), .A1(n4879), .B0(cal_out[361]), .B1(n4908), 
        .Y(n4816) );
  AOI222X1 U9792 ( .A0(cal_out[161]), .A1(n4916), .B0(cal_out[241]), .B1(n4881), .C0(cal_out[201]), .C1(n4912), .Y(n4815) );
  AOI22X1 U9793 ( .A0(cal_out[321]), .A1(n4884), .B0(cal_out[121]), .B1(n4919), 
        .Y(n4814) );
  NAND4BXL U9794 ( .AN(n4817), .B(n4816), .C(n4815), .D(n4814), .Y(
        value_out[1]) );
  AOI22X1 U9795 ( .A0(cal_out[480]), .A1(n4867), .B0(cal_out[280]), .B1(n4866), 
        .Y(n4821) );
  AOI22X1 U9796 ( .A0(cal_out[560]), .A1(n4869), .B0(cal_out[520]), .B1(n4868), 
        .Y(n4820) );
  AOI22X1 U9797 ( .A0(cal_out[0]), .A1(n4871), .B0(cal_out[440]), .B1(n4870), 
        .Y(n4819) );
  AOI22X1 U9798 ( .A0(cal_out[80]), .A1(n4873), .B0(cal_out[40]), .B1(n4872), 
        .Y(n4818) );
  NAND4X1 U9799 ( .A(n4821), .B(n4820), .C(n4819), .D(n4818), .Y(n4825) );
  AOI22X1 U9800 ( .A0(cal_out[400]), .A1(n4879), .B0(cal_out[360]), .B1(n4878), 
        .Y(n4824) );
  AOI222X1 U9801 ( .A0(cal_out[160]), .A1(n4882), .B0(cal_out[240]), .B1(n4881), .C0(cal_out[200]), .C1(n4912), .Y(n4823) );
  AOI22X1 U9802 ( .A0(cal_out[320]), .A1(n4884), .B0(cal_out[120]), .B1(n4883), 
        .Y(n4822) );
  NAND4BXL U9803 ( .AN(n4825), .B(n4824), .C(n4823), .D(n4822), .Y(
        value_out[0]) );
  AOI22X1 U9804 ( .A0(length_reg[77]), .A1(n4867), .B0(length_reg[47]), .B1(
        n4892), .Y(n4829) );
  AOI22X1 U9805 ( .A0(length_reg[89]), .A1(n4869), .B0(length_reg[83]), .B1(
        n4896), .Y(n4828) );
  AOI22X1 U9806 ( .A0(length_reg[5]), .A1(n4871), .B0(length_reg[71]), .B1(
        n4900), .Y(n4827) );
  AOI22X1 U9807 ( .A0(length_reg[17]), .A1(n4873), .B0(length_reg[11]), .B1(
        n4904), .Y(n4826) );
  NAND4X1 U9808 ( .A(n4829), .B(n4828), .C(n4827), .D(n4826), .Y(n4833) );
  AOI22X1 U9809 ( .A0(length_reg[65]), .A1(n4879), .B0(length_reg[59]), .B1(
        n4908), .Y(n4832) );
  AOI222X1 U9810 ( .A0(length_reg[29]), .A1(n4917), .B0(length_reg[41]), .B1(
        n4881), .C0(length_reg[35]), .C1(n4912), .Y(n4831) );
  AOI22X1 U9811 ( .A0(length_reg[53]), .A1(n4884), .B0(length_reg[23]), .B1(
        n4919), .Y(n4830) );
  NAND4BXL U9812 ( .AN(n4833), .B(n4832), .C(n4831), .D(n4830), .Y(
        length_out[5]) );
  AOI22X1 U9813 ( .A0(length_reg[76]), .A1(n4867), .B0(length_reg[46]), .B1(
        n4892), .Y(n4837) );
  AOI22X1 U9814 ( .A0(length_reg[88]), .A1(n4869), .B0(length_reg[82]), .B1(
        n4896), .Y(n4836) );
  AOI22X1 U9815 ( .A0(length_reg[4]), .A1(n4871), .B0(length_reg[70]), .B1(
        n4900), .Y(n4835) );
  AOI22X1 U9816 ( .A0(length_reg[16]), .A1(n4873), .B0(length_reg[10]), .B1(
        n4904), .Y(n4834) );
  NAND4X1 U9817 ( .A(n4837), .B(n4836), .C(n4835), .D(n4834), .Y(n4841) );
  AOI22X1 U9818 ( .A0(length_reg[64]), .A1(n4879), .B0(length_reg[58]), .B1(
        n4908), .Y(n4840) );
  AOI222X1 U9819 ( .A0(length_reg[28]), .A1(n4917), .B0(length_reg[40]), .B1(
        n4881), .C0(length_reg[34]), .C1(n4912), .Y(n4839) );
  AOI22X1 U9820 ( .A0(length_reg[52]), .A1(n4884), .B0(length_reg[22]), .B1(
        n4919), .Y(n4838) );
  NAND4BXL U9821 ( .AN(n4841), .B(n4840), .C(n4839), .D(n4838), .Y(
        length_out[4]) );
  AOI22X1 U9822 ( .A0(length_reg[75]), .A1(n4867), .B0(length_reg[45]), .B1(
        n4866), .Y(n4845) );
  AOI22X1 U9823 ( .A0(length_reg[87]), .A1(n4869), .B0(length_reg[81]), .B1(
        n4868), .Y(n4844) );
  AOI22X1 U9824 ( .A0(length_reg[3]), .A1(n4871), .B0(length_reg[69]), .B1(
        n4870), .Y(n4843) );
  AOI22X1 U9825 ( .A0(length_reg[15]), .A1(n4873), .B0(length_reg[9]), .B1(
        n4872), .Y(n4842) );
  NAND4X1 U9826 ( .A(n4845), .B(n4844), .C(n4843), .D(n4842), .Y(n4849) );
  AOI22X1 U9827 ( .A0(length_reg[63]), .A1(n4879), .B0(length_reg[57]), .B1(
        n4878), .Y(n4848) );
  AOI222X1 U9828 ( .A0(length_reg[27]), .A1(n4917), .B0(length_reg[39]), .B1(
        n4881), .C0(length_reg[33]), .C1(n4912), .Y(n4847) );
  AOI22X1 U9829 ( .A0(length_reg[51]), .A1(n4884), .B0(length_reg[21]), .B1(
        n4883), .Y(n4846) );
  NAND4BXL U9830 ( .AN(n4849), .B(n4848), .C(n4847), .D(n4846), .Y(
        length_out[3]) );
  AOI22X1 U9831 ( .A0(length_reg[74]), .A1(n4867), .B0(length_reg[44]), .B1(
        n4892), .Y(n4853) );
  AOI22X1 U9832 ( .A0(length_reg[86]), .A1(n4869), .B0(length_reg[80]), .B1(
        n4896), .Y(n4852) );
  AOI22X1 U9833 ( .A0(length_reg[2]), .A1(n4871), .B0(length_reg[68]), .B1(
        n4900), .Y(n4851) );
  AOI22X1 U9834 ( .A0(length_reg[14]), .A1(n4873), .B0(length_reg[8]), .B1(
        n4904), .Y(n4850) );
  NAND4X1 U9835 ( .A(n4853), .B(n4852), .C(n4851), .D(n4850), .Y(n4857) );
  AOI22X1 U9836 ( .A0(length_reg[62]), .A1(n4879), .B0(length_reg[56]), .B1(
        n4908), .Y(n4856) );
  AOI222X1 U9837 ( .A0(length_reg[26]), .A1(n4916), .B0(length_reg[38]), .B1(
        n4881), .C0(length_reg[32]), .C1(n4912), .Y(n4855) );
  AOI22X1 U9838 ( .A0(length_reg[50]), .A1(n4884), .B0(length_reg[20]), .B1(
        n4919), .Y(n4854) );
  NAND4BXL U9839 ( .AN(n4857), .B(n4856), .C(n4855), .D(n4854), .Y(
        length_out[2]) );
  AOI22X1 U9840 ( .A0(length_reg[73]), .A1(n4867), .B0(length_reg[43]), .B1(
        n4892), .Y(n4861) );
  AOI22X1 U9841 ( .A0(length_reg[85]), .A1(n4869), .B0(length_reg[79]), .B1(
        n4896), .Y(n4860) );
  AOI22X1 U9842 ( .A0(length_reg[1]), .A1(n4902), .B0(length_reg[67]), .B1(
        n4900), .Y(n4859) );
  AOI22X1 U9843 ( .A0(length_reg[13]), .A1(n4873), .B0(length_reg[7]), .B1(
        n4904), .Y(n4858) );
  NAND4X1 U9844 ( .A(n4861), .B(n4860), .C(n4859), .D(n4858), .Y(n4865) );
  AOI22X1 U9845 ( .A0(length_reg[61]), .A1(n4879), .B0(length_reg[55]), .B1(
        n4908), .Y(n4864) );
  AOI222X1 U9846 ( .A0(length_reg[25]), .A1(n4916), .B0(length_reg[37]), .B1(
        n4881), .C0(length_reg[31]), .C1(n4912), .Y(n4863) );
  AOI22X1 U9847 ( .A0(length_reg[49]), .A1(n4884), .B0(length_reg[19]), .B1(
        n4919), .Y(n4862) );
  NAND4BXL U9848 ( .AN(n4865), .B(n4864), .C(n4863), .D(n4862), .Y(
        length_out[1]) );
  AOI22X1 U9849 ( .A0(length_reg[72]), .A1(n4867), .B0(length_reg[42]), .B1(
        n4892), .Y(n4877) );
  AOI22X1 U9850 ( .A0(length_reg[84]), .A1(n4869), .B0(length_reg[78]), .B1(
        n4896), .Y(n4876) );
  AOI22X1 U9851 ( .A0(length_reg[0]), .A1(n4871), .B0(length_reg[66]), .B1(
        n4900), .Y(n4875) );
  AOI22X1 U9852 ( .A0(length_reg[12]), .A1(n4873), .B0(length_reg[6]), .B1(
        n4904), .Y(n4874) );
  NAND4X1 U9853 ( .A(n4877), .B(n4876), .C(n4875), .D(n4874), .Y(n4888) );
  AOI22X1 U9854 ( .A0(length_reg[60]), .A1(n4879), .B0(length_reg[54]), .B1(
        n4908), .Y(n4887) );
  AOI222X1 U9855 ( .A0(length_reg[24]), .A1(n4916), .B0(length_reg[36]), .B1(
        n4881), .C0(length_reg[30]), .C1(n4912), .Y(n4886) );
  AOI22X1 U9856 ( .A0(length_reg[48]), .A1(n4884), .B0(length_reg[18]), .B1(
        n4919), .Y(n4885) );
  NAND4BXL U9857 ( .AN(n4888), .B(n4887), .C(n4886), .D(n4885), .Y(
        length_out[0]) );
  INVX1 U9858 ( .A(in_cnt_64[0]), .Y(N1034) );
  XOR2X1 U9859 ( .A(add_220_carry[5]), .B(in_cnt_64[5]), .Y(N1039) );
  INVX1 U9860 ( .A(in_matrix_cnt[0]), .Y(N1085) );
  XOR2X1 U9861 ( .A(add_250_carry[4]), .B(N1276), .Y(N1089) );
  NOR2X1 U9862 ( .A(mem_num_0), .B(n5061), .Y(N1233) );
  AOI21X1 U9863 ( .A0(mem_num_0), .A1(n5061), .B0(N1233), .Y(n5639) );
  INVX1 U9864 ( .A(n5639), .Y(N1232) );
  XOR2X1 U9865 ( .A(n5064), .B(N1233), .Y(N1234) );
  INVX1 U9866 ( .A(length_out[0]), .Y(N14358) );
  OAI2BB1X1 U9867 ( .A0N(length_out[0]), .A1N(length_out[1]), .B0(n5640), .Y(
        N14359) );
  OR2X1 U9868 ( .A(n5640), .B(length_out[2]), .Y(n5641) );
  OAI2BB1X1 U9869 ( .A0N(n5640), .A1N(length_out[2]), .B0(n5641), .Y(N14360)
         );
  OR2X1 U9870 ( .A(n5641), .B(length_out[3]), .Y(n5642) );
  OAI2BB1X1 U9871 ( .A0N(n5641), .A1N(length_out[3]), .B0(n5642), .Y(N14361)
         );
  XNOR2X1 U9872 ( .A(length_out[4]), .B(n5642), .Y(N14362) );
  NOR2X1 U9873 ( .A(length_out[4]), .B(n5642), .Y(n5643) );
  XOR2X1 U9874 ( .A(length_out[5]), .B(n5643), .Y(N14363) );
  OAI2BB1X1 U9875 ( .A0N(out_cnt[0]), .A1N(out_cnt[1]), .B0(n5644), .Y(N14365)
         );
  OR2X1 U9876 ( .A(n5644), .B(out_cnt[2]), .Y(n5645) );
  OAI2BB1X1 U9877 ( .A0N(n5644), .A1N(out_cnt[2]), .B0(n5645), .Y(N14366) );
  OR2X1 U9878 ( .A(n5645), .B(out_cnt[3]), .Y(n5646) );
  OAI2BB1X1 U9879 ( .A0N(n5645), .A1N(out_cnt[3]), .B0(n5646), .Y(N14367) );
  XNOR2X1 U9880 ( .A(out_cnt[4]), .B(n5646), .Y(N14368) );
  NOR2X1 U9881 ( .A(out_cnt[4]), .B(n5646), .Y(n5647) );
  XOR2X1 U9882 ( .A(out_cnt[5]), .B(n5647), .Y(N14369) );
  NOR2X1 U9883 ( .A(calin_cnt[4]), .B(calin_cnt[3]), .Y(n5648) );
  OAI21XL U9884 ( .A0(n5064), .A1(n5653), .B0(n5648), .Y(n5649) );
  AOI2BB1X1 U9885 ( .A0N(n5887), .A1N(calin_cnt[1]), .B0(calout_num_0_), .Y(
        n5650) );
  AOI22X1 U9886 ( .A0(calin_cnt[1]), .A1(n5887), .B0(n5650), .B1(calin_cnt[0]), 
        .Y(n5651) );
  AOI32X1 U9887 ( .A0(n5654), .A1(n5653), .A2(n5064), .B0(n5651), .B1(n5654), 
        .Y(n5652) );
  OR4X1 U9888 ( .A(calin_cnt[5]), .B(n5652), .C(calin_cnt[7]), .D(calin_cnt[6]), .Y(r1350_GE_LT_GT_LE) );
  NAND2BX1 U9889 ( .AN(n5086), .B(n5064), .Y(n5655) );
  AOI32X1 U9890 ( .A0(n5087), .A1(n5663), .A2(n5655), .B0(n5887), .B1(n5086), 
        .Y(n5659) );
  OAI21XL U9891 ( .A0(n5087), .A1(n5663), .B0(n5655), .Y(n5658) );
  AOI2BB1X1 U9892 ( .A0N(n5662), .A1N(n5088), .B0(calout_num_0_), .Y(n5656) );
  AOI22X1 U9893 ( .A0(n5088), .A1(n5662), .B0(n5656), .B1(cal_cnt[0]), .Y(
        n5657) );
  AOI22X1 U9894 ( .A0(n5659), .A1(n5658), .B0(n5657), .B1(n5659), .Y(n5661) );
  OR3XL U9895 ( .A(cal_cnt[7]), .B(cal_cnt[6]), .C(cal_cnt[5]), .Y(n5660) );
  OR3XL U9896 ( .A(cal_cnt[4]), .B(n5661), .C(n5660), .Y(N14263) );
endmodule


module MMSA_DW_mult_uns_0 ( a, b, product );
  input [3:0] a;
  input [4:0] b;
  output [8:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n47, n48, n49, n50, n51, n52, n53;

  ADDHXL U2 ( .A(n7), .B(n2), .CO(product[8]), .S(product[7]) );
  ADDFX2 U4 ( .A(n13), .B(n8), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFX2 U5 ( .A(n15), .B(n11), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFX2 U6 ( .A(n14), .B(n9), .CI(n6), .CO(n5), .S(product[3]) );
  ADDHXL U7 ( .A(n12), .B(n16), .CO(n6), .S(product[2]) );
  CMPR22X1 U30 ( .A(n10), .B(n3), .CO(n2), .S(product[6]) );
  INVX1 U31 ( .A(b[0]), .Y(n52) );
  INVX1 U32 ( .A(b[4]), .Y(n53) );
  INVX1 U33 ( .A(b[2]), .Y(n51) );
  INVX1 U34 ( .A(a[1]), .Y(n48) );
  INVX1 U35 ( .A(a[0]), .Y(n47) );
  INVX1 U36 ( .A(a[2]), .Y(n49) );
  INVX1 U37 ( .A(a[3]), .Y(n50) );
  NOR2X1 U38 ( .A(n48), .B(n52), .Y(product[1]) );
  NOR2X1 U39 ( .A(n52), .B(n47), .Y(product[0]) );
  NOR2X1 U40 ( .A(n52), .B(n50), .Y(n9) );
  NOR2X1 U41 ( .A(n50), .B(n51), .Y(n8) );
  NOR2X1 U42 ( .A(n50), .B(n53), .Y(n7) );
  NOR2X1 U43 ( .A(n47), .B(n51), .Y(n16) );
  NOR2X1 U44 ( .A(n47), .B(n53), .Y(n15) );
  NOR2X1 U45 ( .A(n48), .B(n51), .Y(n14) );
  NOR2X1 U46 ( .A(n48), .B(n53), .Y(n13) );
  NOR2X1 U47 ( .A(n52), .B(n49), .Y(n12) );
  NOR2X1 U48 ( .A(n51), .B(n49), .Y(n11) );
  NOR2X1 U49 ( .A(n53), .B(n49), .Y(n10) );
endmodule


module MMSA_DW_mult_uns_1 ( a, b, product );
  input [3:0] a;
  input [4:0] b;
  output [8:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n47, n48, n49, n50, n51, n52, n53;

  ADDHXL U2 ( .A(n7), .B(n2), .CO(product[8]), .S(product[7]) );
  ADDFX2 U4 ( .A(n13), .B(n8), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFX2 U5 ( .A(n15), .B(n11), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFX2 U6 ( .A(n14), .B(n9), .CI(n6), .CO(n5), .S(product[3]) );
  ADDHXL U7 ( .A(n12), .B(n16), .CO(n6), .S(product[2]) );
  CMPR22X1 U30 ( .A(n10), .B(n3), .CO(n2), .S(product[6]) );
  INVX1 U31 ( .A(b[0]), .Y(n52) );
  INVX1 U32 ( .A(b[4]), .Y(n53) );
  INVX1 U33 ( .A(b[2]), .Y(n51) );
  INVX1 U34 ( .A(a[1]), .Y(n48) );
  INVX1 U35 ( .A(a[0]), .Y(n47) );
  INVX1 U36 ( .A(a[2]), .Y(n49) );
  INVX1 U37 ( .A(a[3]), .Y(n50) );
  NOR2X1 U38 ( .A(n48), .B(n52), .Y(product[1]) );
  NOR2X1 U39 ( .A(n52), .B(n47), .Y(product[0]) );
  NOR2X1 U40 ( .A(n52), .B(n50), .Y(n9) );
  NOR2X1 U41 ( .A(n50), .B(n51), .Y(n8) );
  NOR2X1 U42 ( .A(n50), .B(n53), .Y(n7) );
  NOR2X1 U43 ( .A(n47), .B(n51), .Y(n16) );
  NOR2X1 U44 ( .A(n47), .B(n53), .Y(n15) );
  NOR2X1 U45 ( .A(n48), .B(n51), .Y(n14) );
  NOR2X1 U46 ( .A(n48), .B(n53), .Y(n13) );
  NOR2X1 U47 ( .A(n52), .B(n49), .Y(n12) );
  NOR2X1 U48 ( .A(n51), .B(n49), .Y(n11) );
  NOR2X1 U49 ( .A(n53), .B(n49), .Y(n10) );
endmodule


module MMSA_DW01_add_8 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_add_9 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NOR2X1 U2 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U3 ( .A(B[0]), .Y(n2) );
  INVX1 U4 ( .A(A[0]), .Y(n1) );
endmodule


module MMSA_DW01_add_10 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NOR2X1 U2 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U3 ( .A(B[0]), .Y(n2) );
  INVX1 U4 ( .A(A[0]), .Y(n1) );
endmodule


module MMSA_DW01_add_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_add_2 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_add_3 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NOR2X1 U2 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U3 ( .A(B[0]), .Y(n2) );
  INVX1 U4 ( .A(A[0]), .Y(n1) );
endmodule


module MMSA_DW01_add_4 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_add_5 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_add_6 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_add_7 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_6 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  CMPR22X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CMPR22X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_4 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  CMPR22X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  CMPR22X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CMPR22X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_3 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  CMPR22X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  CMPR22X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CMPR22X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_2 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  CMPR22X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  CMPR22X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CMPR22X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CMPR22X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CMPR22X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CMPR22X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_1 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_1_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_1_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_1_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_2 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_2_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_2_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_2_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_3 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_3_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_3_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_3_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_4 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_4_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_4_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_4_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_5 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_5_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_5_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_5_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_6 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_6_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_6_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_6_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_6_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_7 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_7_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_7_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_7_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_7_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_8 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_8_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_8_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_8_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_8_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n658), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n657), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n656), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n661), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n662), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n660), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n659), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n659) );
  INVX1 U492 ( .A(n121), .Y(n662) );
  INVX1 U493 ( .A(n96), .Y(n656) );
  INVX1 U494 ( .A(n82), .Y(n658) );
  INVX1 U495 ( .A(n648), .Y(n679) );
  CLKINVX3 U496 ( .A(n709), .Y(n678) );
  CLKINVX3 U497 ( .A(n651), .Y(n670) );
  CLKINVX3 U498 ( .A(n649), .Y(n676) );
  CLKINVX3 U499 ( .A(n650), .Y(n673) );
  CLKINVX3 U500 ( .A(n647), .Y(n663) );
  CLKINVX3 U501 ( .A(n652), .Y(n667) );
  CLKINVX3 U502 ( .A(n653), .Y(n686) );
  CLKINVX3 U503 ( .A(n654), .Y(n684) );
  INVX1 U504 ( .A(n655), .Y(n681) );
  INVX1 U505 ( .A(n728), .Y(n674) );
  INVX1 U506 ( .A(n710), .Y(n677) );
  INVX1 U507 ( .A(n712), .Y(n675) );
  INVX1 U508 ( .A(n730), .Y(n672) );
  INVX1 U509 ( .A(n140), .Y(n660) );
  INVX1 U510 ( .A(n764), .Y(n668) );
  INVX1 U511 ( .A(n746), .Y(n671) );
  INVX1 U512 ( .A(n748), .Y(n669) );
  INVX1 U513 ( .A(n108), .Y(n661) );
  INVX1 U514 ( .A(n782), .Y(n666) );
  INVX1 U515 ( .A(n766), .Y(n664) );
  INVX1 U516 ( .A(n784), .Y(n665) );
  INVX1 U517 ( .A(n798), .Y(n685) );
  INVX1 U518 ( .A(n88), .Y(n657) );
  INVX1 U519 ( .A(n814), .Y(n682) );
  INVX1 U520 ( .A(n800), .Y(n683) );
  INVX1 U521 ( .A(n816), .Y(n680) );
  XOR2X2 U522 ( .A(a[2]), .B(n679), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n673), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n676), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n670), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n687) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n667), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n686), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n684), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n687), .B(n663), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n665), .B0(n666), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n683), .B0(n685), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n680), .B0(n682), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n678), .B0(n694), .B1(n687), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n678), .B0(n695), .B1(n687), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n678), .B0(n696), .B1(n687), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n678), .B0(n697), .B1(n687), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n678), .B0(n698), .B1(n687), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n678), .B0(n699), .B1(n687), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n678), .B0(n700), .B1(n687), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n678), .B0(n701), .B1(n687), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n678), .B0(n702), .B1(n687), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n678), .B0(n703), .B1(n687), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n678), .B0(n704), .B1(n687), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n678), .B0(n705), .B1(n687), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n678), .B0(n706), .B1(n687), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n678), .B0(n707), .B1(n687), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n678), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n679), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n663), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n677), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n677), .B0(n675), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n663), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n674), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n674), .B0(n672), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n663), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n671), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n671), .B0(n669), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n670), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n663), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n668), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n668), .B0(n664), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n663), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n666), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n666), .B0(n665), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n686), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n663), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n685), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n685), .B0(n683), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n684), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n663), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n682), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n682), .B0(n680), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n681), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n679), .B0(n678), .Y(n267) );
  NOR2X1 U793 ( .A(n679), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n676), .A1(n647), .A2(n710), .B0(n676), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n673), .A1(n647), .A2(n728), .B0(n673), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n670), .A1(n647), .A2(n746), .B0(n670), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n667), .A1(n647), .A2(n764), .B0(n667), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n686), .A1(n647), .A2(n782), .B0(n686), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n684), .A1(n647), .A2(n798), .B0(n684), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n681), .A1(n647), .A2(n814), .B0(n681), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n681), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n670), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n684), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n675), .B0(n677), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n676), .Y(n727) );
  XNOR2X1 U814 ( .A(n676), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n672), .B0(n674), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n673), .Y(n745) );
  XNOR2X1 U818 ( .A(n673), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n686), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n664), .B0(n668), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n667), .Y(n781) );
  XNOR2X1 U826 ( .A(n667), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_9 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_9_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_9_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_9_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_9_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_10 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_10_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_10_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_10_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_10_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_11 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_11_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_11_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_11_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_11_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_12 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_12_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_12_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_12_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_12_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_13 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_13_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_13_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_13_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_13_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_14 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_14_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_14_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_14_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_14_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_15 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_15_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_15_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_15_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_15_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_16 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_16_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_16_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_16_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_16_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n658), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n657), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n656), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n661), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n662), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n660), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n659), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n659) );
  INVX1 U492 ( .A(n121), .Y(n662) );
  INVX1 U493 ( .A(n96), .Y(n656) );
  INVX1 U494 ( .A(n82), .Y(n658) );
  INVX1 U495 ( .A(n648), .Y(n686) );
  CLKINVX3 U496 ( .A(n709), .Y(n685) );
  CLKINVX3 U497 ( .A(n651), .Y(n677) );
  CLKINVX3 U498 ( .A(n649), .Y(n683) );
  CLKINVX3 U499 ( .A(n650), .Y(n680) );
  CLKINVX3 U500 ( .A(n647), .Y(n663) );
  CLKINVX3 U501 ( .A(n652), .Y(n674) );
  CLKINVX3 U502 ( .A(n653), .Y(n671) );
  CLKINVX3 U503 ( .A(n654), .Y(n668) );
  INVX1 U504 ( .A(n655), .Y(n665) );
  INVX1 U505 ( .A(n728), .Y(n681) );
  INVX1 U506 ( .A(n710), .Y(n684) );
  INVX1 U507 ( .A(n712), .Y(n682) );
  INVX1 U508 ( .A(n730), .Y(n679) );
  INVX1 U509 ( .A(n140), .Y(n660) );
  INVX1 U510 ( .A(n764), .Y(n675) );
  INVX1 U511 ( .A(n746), .Y(n678) );
  INVX1 U512 ( .A(n748), .Y(n676) );
  INVX1 U513 ( .A(n108), .Y(n661) );
  INVX1 U514 ( .A(n782), .Y(n672) );
  INVX1 U515 ( .A(n766), .Y(n673) );
  INVX1 U516 ( .A(n784), .Y(n670) );
  INVX1 U517 ( .A(n798), .Y(n669) );
  INVX1 U518 ( .A(n88), .Y(n657) );
  INVX1 U519 ( .A(n814), .Y(n666) );
  INVX1 U520 ( .A(n800), .Y(n667) );
  INVX1 U521 ( .A(n816), .Y(n664) );
  XOR2X2 U522 ( .A(a[2]), .B(n686), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n680), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n683), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n677), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n687) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n674), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n671), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n668), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n687), .B(n663), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n670), .B0(n672), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n667), .B0(n669), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n664), .B0(n666), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n685), .B0(n694), .B1(n687), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n685), .B0(n695), .B1(n687), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n685), .B0(n696), .B1(n687), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n685), .B0(n697), .B1(n687), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n685), .B0(n698), .B1(n687), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n685), .B0(n699), .B1(n687), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n685), .B0(n700), .B1(n687), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n685), .B0(n701), .B1(n687), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n685), .B0(n702), .B1(n687), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n685), .B0(n703), .B1(n687), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n685), .B0(n704), .B1(n687), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n685), .B0(n705), .B1(n687), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n685), .B0(n706), .B1(n687), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n685), .B0(n707), .B1(n687), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n685), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n686), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n663), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n684), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n684), .B0(n682), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n663), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n681), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n681), .B0(n679), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n663), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n678), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n678), .B0(n676), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n677), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n663), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n675), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n675), .B0(n673), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n663), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n672), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n672), .B0(n670), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n671), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n663), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n669), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n669), .B0(n667), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n668), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n663), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n666), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n666), .B0(n664), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n665), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n686), .B0(n685), .Y(n267) );
  NOR2X1 U793 ( .A(n686), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n683), .A1(n647), .A2(n710), .B0(n683), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n680), .A1(n647), .A2(n728), .B0(n680), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n677), .A1(n647), .A2(n746), .B0(n677), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n674), .A1(n647), .A2(n764), .B0(n674), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n671), .A1(n647), .A2(n782), .B0(n671), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n668), .A1(n647), .A2(n798), .B0(n668), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n665), .A1(n647), .A2(n814), .B0(n665), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n665), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n677), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n668), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n682), .B0(n684), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n683), .Y(n727) );
  XNOR2X1 U814 ( .A(n683), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n679), .B0(n681), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n680), .Y(n745) );
  XNOR2X1 U818 ( .A(n680), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n671), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n673), .B0(n675), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n674), .Y(n781) );
  XNOR2X1 U826 ( .A(n674), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_17 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_17_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_17_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_17_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_17_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_18 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_18_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_18_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_18_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_18_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_19 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_19_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_19_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_19_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_19_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_20 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_20_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_20_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_20_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_20_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_21 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_21_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_21_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_21_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_21_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_22 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_22_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_22_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_22_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_22_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_23 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_23_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_23_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_23_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_23_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_24 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_24_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_24_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_24_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_24_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n658), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n657), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n656), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n661), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n662), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n660), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n659), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n659) );
  INVX1 U492 ( .A(n121), .Y(n662) );
  INVX1 U493 ( .A(n96), .Y(n656) );
  INVX1 U494 ( .A(n82), .Y(n658) );
  INVX1 U495 ( .A(n648), .Y(n686) );
  CLKINVX3 U496 ( .A(n709), .Y(n685) );
  CLKINVX3 U497 ( .A(n651), .Y(n677) );
  CLKINVX3 U498 ( .A(n649), .Y(n683) );
  CLKINVX3 U499 ( .A(n650), .Y(n680) );
  CLKINVX3 U500 ( .A(n647), .Y(n663) );
  CLKINVX3 U501 ( .A(n652), .Y(n674) );
  CLKINVX3 U502 ( .A(n653), .Y(n671) );
  CLKINVX3 U503 ( .A(n654), .Y(n668) );
  INVX1 U504 ( .A(n655), .Y(n665) );
  INVX1 U505 ( .A(n728), .Y(n681) );
  INVX1 U506 ( .A(n710), .Y(n684) );
  INVX1 U507 ( .A(n712), .Y(n682) );
  INVX1 U508 ( .A(n730), .Y(n679) );
  INVX1 U509 ( .A(n140), .Y(n660) );
  INVX1 U510 ( .A(n764), .Y(n675) );
  INVX1 U511 ( .A(n746), .Y(n678) );
  INVX1 U512 ( .A(n748), .Y(n676) );
  INVX1 U513 ( .A(n108), .Y(n661) );
  INVX1 U514 ( .A(n782), .Y(n672) );
  INVX1 U515 ( .A(n766), .Y(n673) );
  INVX1 U516 ( .A(n784), .Y(n670) );
  INVX1 U517 ( .A(n798), .Y(n669) );
  INVX1 U518 ( .A(n88), .Y(n657) );
  INVX1 U519 ( .A(n814), .Y(n666) );
  INVX1 U520 ( .A(n800), .Y(n667) );
  INVX1 U521 ( .A(n816), .Y(n664) );
  XOR2X2 U522 ( .A(a[2]), .B(n686), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n680), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n683), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n677), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n687) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n674), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n671), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n668), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n687), .B(n663), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n670), .B0(n672), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n667), .B0(n669), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n664), .B0(n666), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n685), .B0(n694), .B1(n687), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n685), .B0(n695), .B1(n687), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n685), .B0(n696), .B1(n687), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n685), .B0(n697), .B1(n687), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n685), .B0(n698), .B1(n687), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n685), .B0(n699), .B1(n687), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n685), .B0(n700), .B1(n687), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n685), .B0(n701), .B1(n687), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n685), .B0(n702), .B1(n687), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n685), .B0(n703), .B1(n687), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n685), .B0(n704), .B1(n687), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n685), .B0(n705), .B1(n687), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n685), .B0(n706), .B1(n687), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n685), .B0(n707), .B1(n687), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n685), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n686), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n663), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n684), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n684), .B0(n682), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n663), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n681), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n681), .B0(n679), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n663), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n678), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n678), .B0(n676), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n677), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n663), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n675), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n675), .B0(n673), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n663), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n672), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n672), .B0(n670), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n671), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n663), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n669), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n669), .B0(n667), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n668), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n663), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n666), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n666), .B0(n664), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n665), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n686), .B0(n685), .Y(n267) );
  NOR2X1 U793 ( .A(n686), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n683), .A1(n647), .A2(n710), .B0(n683), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n680), .A1(n647), .A2(n728), .B0(n680), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n677), .A1(n647), .A2(n746), .B0(n677), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n674), .A1(n647), .A2(n764), .B0(n674), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n671), .A1(n647), .A2(n782), .B0(n671), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n668), .A1(n647), .A2(n798), .B0(n668), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n665), .A1(n647), .A2(n814), .B0(n665), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n665), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n677), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n668), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n682), .B0(n684), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n683), .Y(n727) );
  XNOR2X1 U814 ( .A(n683), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n679), .B0(n681), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n680), .Y(n745) );
  XNOR2X1 U818 ( .A(n680), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n671), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n673), .B0(n675), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n674), .Y(n781) );
  XNOR2X1 U826 ( .A(n674), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_25 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_25_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_25_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_25_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_25_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_26 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_26_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_26_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_26_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_26_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_27 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_27_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_27_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_27_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_27_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_28 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_28_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_28_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_28_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_28_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_29 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_29_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_29_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_29_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_29_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_30 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_30_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_30_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_30_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_30_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_31 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_31_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_31_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_31_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_31_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_32 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_32_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_32_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_32_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n658), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n657), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n656), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n661), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n662), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n660), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n659), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n659) );
  INVX1 U492 ( .A(n121), .Y(n662) );
  INVX1 U493 ( .A(n96), .Y(n656) );
  INVX1 U494 ( .A(n82), .Y(n658) );
  INVX1 U495 ( .A(n648), .Y(n686) );
  CLKINVX3 U496 ( .A(n709), .Y(n685) );
  CLKINVX3 U497 ( .A(n651), .Y(n677) );
  CLKINVX3 U498 ( .A(n649), .Y(n683) );
  CLKINVX3 U499 ( .A(n650), .Y(n680) );
  CLKINVX3 U500 ( .A(n647), .Y(n663) );
  CLKINVX3 U501 ( .A(n652), .Y(n674) );
  CLKINVX3 U502 ( .A(n653), .Y(n671) );
  CLKINVX3 U503 ( .A(n654), .Y(n668) );
  INVX1 U504 ( .A(n655), .Y(n665) );
  INVX1 U505 ( .A(n728), .Y(n681) );
  INVX1 U506 ( .A(n710), .Y(n684) );
  INVX1 U507 ( .A(n712), .Y(n682) );
  INVX1 U508 ( .A(n730), .Y(n679) );
  INVX1 U509 ( .A(n140), .Y(n660) );
  INVX1 U510 ( .A(n764), .Y(n675) );
  INVX1 U511 ( .A(n746), .Y(n678) );
  INVX1 U512 ( .A(n748), .Y(n676) );
  INVX1 U513 ( .A(n108), .Y(n661) );
  INVX1 U514 ( .A(n782), .Y(n672) );
  INVX1 U515 ( .A(n766), .Y(n673) );
  INVX1 U516 ( .A(n784), .Y(n670) );
  INVX1 U517 ( .A(n798), .Y(n669) );
  INVX1 U518 ( .A(n88), .Y(n657) );
  INVX1 U519 ( .A(n814), .Y(n666) );
  INVX1 U520 ( .A(n800), .Y(n667) );
  INVX1 U521 ( .A(n816), .Y(n664) );
  XOR2X2 U522 ( .A(a[2]), .B(n686), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n680), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n683), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n677), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n687) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n674), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n671), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n668), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n687), .B(n663), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n670), .B0(n672), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n667), .B0(n669), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n664), .B0(n666), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n685), .B0(n694), .B1(n687), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n685), .B0(n695), .B1(n687), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n685), .B0(n696), .B1(n687), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n685), .B0(n697), .B1(n687), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n685), .B0(n698), .B1(n687), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n685), .B0(n699), .B1(n687), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n685), .B0(n700), .B1(n687), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n685), .B0(n701), .B1(n687), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n685), .B0(n702), .B1(n687), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n685), .B0(n703), .B1(n687), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n685), .B0(n704), .B1(n687), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n685), .B0(n705), .B1(n687), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n685), .B0(n706), .B1(n687), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n685), .B0(n707), .B1(n687), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n685), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n686), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n663), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n684), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n684), .B0(n682), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n663), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n681), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n681), .B0(n679), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n663), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n678), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n678), .B0(n676), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n677), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n663), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n675), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n675), .B0(n673), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n663), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n672), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n672), .B0(n670), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n671), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n663), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n669), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n669), .B0(n667), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n668), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n663), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n666), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n666), .B0(n664), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n665), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n686), .B0(n685), .Y(n267) );
  NOR2X1 U793 ( .A(n686), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n683), .A1(n647), .A2(n710), .B0(n683), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n680), .A1(n647), .A2(n728), .B0(n680), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n677), .A1(n647), .A2(n746), .B0(n677), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n674), .A1(n647), .A2(n764), .B0(n674), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n671), .A1(n647), .A2(n782), .B0(n671), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n668), .A1(n647), .A2(n798), .B0(n668), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n665), .A1(n647), .A2(n814), .B0(n665), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n665), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n677), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n668), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n682), .B0(n684), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n683), .Y(n727) );
  XNOR2X1 U814 ( .A(n683), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n679), .B0(n681), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n680), .Y(n745) );
  XNOR2X1 U818 ( .A(n680), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n671), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n673), .B0(n675), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n674), .Y(n781) );
  XNOR2X1 U826 ( .A(n674), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_33 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_33_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_33_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_33_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_33_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_34 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_34_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_34_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_34_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_34_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_35 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_35_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_35_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_35_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_35_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_36 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_36_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_36_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_36_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_36_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_37 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_37_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_37_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_37_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_37_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_38 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_38_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_38_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_38_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_38_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_39 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_39_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_39_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_39_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_39_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_40 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_40_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_40_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_40_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_40_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n658), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n657), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n656), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n661), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n662), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n660), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n659), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n659) );
  INVX1 U492 ( .A(n121), .Y(n662) );
  INVX1 U493 ( .A(n96), .Y(n656) );
  INVX1 U494 ( .A(n82), .Y(n658) );
  INVX1 U495 ( .A(n648), .Y(n679) );
  CLKINVX3 U496 ( .A(n709), .Y(n678) );
  CLKINVX3 U497 ( .A(n651), .Y(n670) );
  CLKINVX3 U498 ( .A(n649), .Y(n676) );
  CLKINVX3 U499 ( .A(n650), .Y(n673) );
  CLKINVX3 U500 ( .A(n647), .Y(n663) );
  CLKINVX3 U501 ( .A(n652), .Y(n667) );
  CLKINVX3 U502 ( .A(n653), .Y(n686) );
  CLKINVX3 U503 ( .A(n654), .Y(n684) );
  INVX1 U504 ( .A(n655), .Y(n681) );
  INVX1 U505 ( .A(n728), .Y(n674) );
  INVX1 U506 ( .A(n710), .Y(n677) );
  INVX1 U507 ( .A(n712), .Y(n675) );
  INVX1 U508 ( .A(n730), .Y(n672) );
  INVX1 U509 ( .A(n140), .Y(n660) );
  INVX1 U510 ( .A(n764), .Y(n668) );
  INVX1 U511 ( .A(n746), .Y(n671) );
  INVX1 U512 ( .A(n748), .Y(n669) );
  INVX1 U513 ( .A(n108), .Y(n661) );
  INVX1 U514 ( .A(n782), .Y(n666) );
  INVX1 U515 ( .A(n766), .Y(n664) );
  INVX1 U516 ( .A(n784), .Y(n665) );
  INVX1 U517 ( .A(n798), .Y(n685) );
  INVX1 U518 ( .A(n88), .Y(n657) );
  INVX1 U519 ( .A(n814), .Y(n682) );
  INVX1 U520 ( .A(n800), .Y(n683) );
  INVX1 U521 ( .A(n816), .Y(n680) );
  XOR2X2 U522 ( .A(a[2]), .B(n679), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n673), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n676), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n670), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n687) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n667), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n686), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n684), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n687), .B(n663), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n665), .B0(n666), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n683), .B0(n685), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n680), .B0(n682), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n678), .B0(n694), .B1(n687), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n678), .B0(n695), .B1(n687), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n678), .B0(n696), .B1(n687), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n678), .B0(n697), .B1(n687), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n678), .B0(n698), .B1(n687), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n678), .B0(n699), .B1(n687), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n678), .B0(n700), .B1(n687), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n678), .B0(n701), .B1(n687), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n678), .B0(n702), .B1(n687), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n678), .B0(n703), .B1(n687), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n678), .B0(n704), .B1(n687), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n678), .B0(n705), .B1(n687), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n678), .B0(n706), .B1(n687), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n678), .B0(n707), .B1(n687), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n678), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n679), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n663), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n677), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n677), .B0(n675), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n663), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n674), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n674), .B0(n672), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n663), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n671), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n671), .B0(n669), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n670), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n663), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n668), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n668), .B0(n664), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n663), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n666), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n666), .B0(n665), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n686), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n663), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n685), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n685), .B0(n683), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n684), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n663), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n682), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n682), .B0(n680), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n681), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n679), .B0(n678), .Y(n267) );
  NOR2X1 U793 ( .A(n679), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n676), .A1(n647), .A2(n710), .B0(n676), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n673), .A1(n647), .A2(n728), .B0(n673), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n670), .A1(n647), .A2(n746), .B0(n670), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n667), .A1(n647), .A2(n764), .B0(n667), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n686), .A1(n647), .A2(n782), .B0(n686), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n684), .A1(n647), .A2(n798), .B0(n684), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n681), .A1(n647), .A2(n814), .B0(n681), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n681), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n670), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n684), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n675), .B0(n677), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n676), .Y(n727) );
  XNOR2X1 U814 ( .A(n676), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n672), .B0(n674), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n673), .Y(n745) );
  XNOR2X1 U818 ( .A(n673), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n686), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n664), .B0(n668), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n667), .Y(n781) );
  XNOR2X1 U826 ( .A(n667), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_41 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_41_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_41_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_41_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_41_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_42 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_42_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_42_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_42_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_42_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_43 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_43_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_43_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_43_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_43_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_44 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_44_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_44_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_44_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_44_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_45 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_45_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_45_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_45_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_45_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_46 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_46_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_46_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_46_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_46_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_47 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_47_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_47_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_47_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_47_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_48 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_48_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_48_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_48_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_48_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n658), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n657), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n656), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n661), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n662), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n660), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n659), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n659) );
  INVX1 U492 ( .A(n121), .Y(n662) );
  INVX1 U493 ( .A(n96), .Y(n656) );
  INVX1 U494 ( .A(n82), .Y(n658) );
  INVX1 U495 ( .A(n648), .Y(n686) );
  CLKINVX3 U496 ( .A(n709), .Y(n685) );
  CLKINVX3 U497 ( .A(n651), .Y(n677) );
  CLKINVX3 U498 ( .A(n649), .Y(n683) );
  CLKINVX3 U499 ( .A(n650), .Y(n680) );
  CLKINVX3 U500 ( .A(n647), .Y(n663) );
  CLKINVX3 U501 ( .A(n652), .Y(n674) );
  CLKINVX3 U502 ( .A(n653), .Y(n671) );
  CLKINVX3 U503 ( .A(n654), .Y(n668) );
  INVX1 U504 ( .A(n655), .Y(n665) );
  INVX1 U505 ( .A(n728), .Y(n681) );
  INVX1 U506 ( .A(n710), .Y(n684) );
  INVX1 U507 ( .A(n712), .Y(n682) );
  INVX1 U508 ( .A(n730), .Y(n679) );
  INVX1 U509 ( .A(n140), .Y(n660) );
  INVX1 U510 ( .A(n764), .Y(n675) );
  INVX1 U511 ( .A(n746), .Y(n678) );
  INVX1 U512 ( .A(n748), .Y(n676) );
  INVX1 U513 ( .A(n108), .Y(n661) );
  INVX1 U514 ( .A(n782), .Y(n672) );
  INVX1 U515 ( .A(n766), .Y(n673) );
  INVX1 U516 ( .A(n784), .Y(n670) );
  INVX1 U517 ( .A(n798), .Y(n669) );
  INVX1 U518 ( .A(n88), .Y(n657) );
  INVX1 U519 ( .A(n814), .Y(n666) );
  INVX1 U520 ( .A(n800), .Y(n667) );
  INVX1 U521 ( .A(n816), .Y(n664) );
  XOR2X2 U522 ( .A(a[2]), .B(n686), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n680), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n683), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n677), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n687) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n674), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n671), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n668), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n687), .B(n663), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n670), .B0(n672), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n667), .B0(n669), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n664), .B0(n666), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n685), .B0(n694), .B1(n687), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n685), .B0(n695), .B1(n687), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n685), .B0(n696), .B1(n687), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n685), .B0(n697), .B1(n687), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n685), .B0(n698), .B1(n687), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n685), .B0(n699), .B1(n687), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n685), .B0(n700), .B1(n687), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n685), .B0(n701), .B1(n687), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n685), .B0(n702), .B1(n687), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n685), .B0(n703), .B1(n687), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n685), .B0(n704), .B1(n687), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n685), .B0(n705), .B1(n687), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n685), .B0(n706), .B1(n687), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n685), .B0(n707), .B1(n687), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n685), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n686), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n663), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n684), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n684), .B0(n682), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n663), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n681), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n681), .B0(n679), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n663), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n678), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n678), .B0(n676), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n677), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n663), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n675), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n675), .B0(n673), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n663), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n672), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n672), .B0(n670), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n671), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n663), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n669), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n669), .B0(n667), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n668), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n663), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n666), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n666), .B0(n664), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n665), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n686), .B0(n685), .Y(n267) );
  NOR2X1 U793 ( .A(n686), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n683), .A1(n647), .A2(n710), .B0(n683), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n680), .A1(n647), .A2(n728), .B0(n680), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n677), .A1(n647), .A2(n746), .B0(n677), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n674), .A1(n647), .A2(n764), .B0(n674), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n671), .A1(n647), .A2(n782), .B0(n671), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n668), .A1(n647), .A2(n798), .B0(n668), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n665), .A1(n647), .A2(n814), .B0(n665), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n665), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n677), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n668), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n682), .B0(n684), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n683), .Y(n727) );
  XNOR2X1 U814 ( .A(n683), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n679), .B0(n681), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n680), .Y(n745) );
  XNOR2X1 U818 ( .A(n680), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n671), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n673), .B0(n675), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n674), .Y(n781) );
  XNOR2X1 U826 ( .A(n674), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_49 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_49_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_49_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_49_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_49_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_50 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_50_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_50_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_50_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_50_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_51 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_51_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_51_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_51_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_51_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_52 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_52_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_52_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_52_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_52_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_53 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_53_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_53_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_53_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_53_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_54 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_54_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_54_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_54_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_54_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  INVX1 U495 ( .A(n648), .Y(n685) );
  CLKINVX3 U496 ( .A(n709), .Y(n684) );
  CLKINVX3 U497 ( .A(n651), .Y(n674) );
  CLKINVX3 U498 ( .A(n649), .Y(n682) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n647), .Y(n687) );
  CLKINVX3 U501 ( .A(n652), .Y(n671) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n655), .Y(n658) );
  INVX1 U505 ( .A(n728), .Y(n679) );
  INVX1 U506 ( .A(n710), .Y(n683) );
  INVX1 U507 ( .A(n712), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n764), .Y(n672) );
  INVX1 U511 ( .A(n746), .Y(n675) );
  INVX1 U512 ( .A(n748), .Y(n673) );
  INVX1 U513 ( .A(n108), .Y(n669) );
  INVX1 U514 ( .A(n782), .Y(n668) );
  INVX1 U515 ( .A(n766), .Y(n670) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n88), .Y(n660) );
  INVX1 U519 ( .A(n814), .Y(n659) );
  INVX1 U520 ( .A(n800), .Y(n661) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n686) );
  BUFX3 U528 ( .A(a[7]), .Y(n651) );
  BUFX3 U529 ( .A(a[3]), .Y(n649) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(b[0]), .Y(n647) );
  XOR2X2 U532 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_55 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_55_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_55_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_55_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_55_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837;

  ADDFX2 U52 ( .A(n268), .B(n655), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n659), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n663), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n668), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n664), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n675), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n679), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n679) );
  INVX1 U492 ( .A(n121), .Y(n664) );
  INVX1 U493 ( .A(n96), .Y(n663) );
  INVX1 U494 ( .A(n82), .Y(n655) );
  INVX1 U495 ( .A(n647), .Y(n684) );
  CLKINVX3 U496 ( .A(n708), .Y(n683) );
  CLKINVX3 U497 ( .A(n650), .Y(n673) );
  CLKINVX3 U498 ( .A(n648), .Y(n681) );
  CLKINVX3 U499 ( .A(n649), .Y(n677) );
  CLKINVX3 U500 ( .A(n651), .Y(n670) );
  CLKINVX3 U501 ( .A(n652), .Y(n666) );
  CLKINVX3 U502 ( .A(n653), .Y(n661) );
  INVX1 U503 ( .A(n654), .Y(n657) );
  INVX1 U504 ( .A(n727), .Y(n678) );
  INVX1 U505 ( .A(n709), .Y(n682) );
  INVX1 U506 ( .A(n711), .Y(n680) );
  INVX1 U507 ( .A(n729), .Y(n676) );
  INVX1 U508 ( .A(n140), .Y(n675) );
  INVX1 U509 ( .A(n763), .Y(n671) );
  INVX1 U510 ( .A(n745), .Y(n674) );
  INVX1 U511 ( .A(n747), .Y(n672) );
  INVX1 U512 ( .A(n108), .Y(n668) );
  INVX1 U513 ( .A(n781), .Y(n667) );
  INVX1 U514 ( .A(n765), .Y(n669) );
  INVX1 U515 ( .A(n783), .Y(n665) );
  INVX1 U516 ( .A(n797), .Y(n662) );
  INVX1 U517 ( .A(n88), .Y(n659) );
  INVX1 U518 ( .A(n813), .Y(n658) );
  INVX1 U519 ( .A(n799), .Y(n660) );
  INVX1 U520 ( .A(n815), .Y(n656) );
  XOR2X2 U521 ( .A(a[2]), .B(n684), .Y(n709) );
  BUFX3 U522 ( .A(a[1]), .Y(n647) );
  XOR2X2 U523 ( .A(a[6]), .B(n677), .Y(n745) );
  XOR2X2 U524 ( .A(a[4]), .B(n681), .Y(n727) );
  XOR2X2 U525 ( .A(a[8]), .B(n673), .Y(n763) );
  CLKINVX3 U526 ( .A(b[0]), .Y(n686) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n685) );
  BUFX3 U528 ( .A(a[7]), .Y(n650) );
  BUFX3 U529 ( .A(a[3]), .Y(n648) );
  BUFX3 U530 ( .A(a[5]), .Y(n649) );
  XOR2X2 U531 ( .A(a[10]), .B(n670), .Y(n781) );
  XOR2X2 U532 ( .A(a[12]), .B(n666), .Y(n797) );
  BUFX3 U533 ( .A(a[9]), .Y(n651) );
  BUFX3 U534 ( .A(a[11]), .Y(n652) );
  BUFX3 U535 ( .A(a[13]), .Y(n653) );
  XOR2X2 U536 ( .A(a[14]), .B(n661), .Y(n813) );
  BUFX3 U537 ( .A(a[15]), .Y(n654) );
  NAND2X4 U538 ( .A(n813), .B(n829), .Y(n815) );
  NAND2X4 U539 ( .A(n745), .B(n832), .Y(n747) );
  NAND2X4 U540 ( .A(n797), .B(n833), .Y(n799) );
  NAND2X4 U541 ( .A(n709), .B(n834), .Y(n711) );
  NAND2X4 U542 ( .A(n727), .B(n835), .Y(n729) );
  NAND2X4 U543 ( .A(n781), .B(n836), .Y(n783) );
  NAND2X4 U544 ( .A(n763), .B(n837), .Y(n765) );
  INVX1 U545 ( .A(n51), .Y(product[31]) );
  NOR2X1 U546 ( .A(n685), .B(n686), .Y(product[0]) );
  AOI22X1 U547 ( .A0(n687), .A1(n665), .B0(n667), .B1(n688), .Y(n96) );
  AOI22X1 U548 ( .A0(n689), .A1(n660), .B0(n662), .B1(n690), .Y(n88) );
  AOI22X1 U549 ( .A0(n691), .A1(n656), .B0(n658), .B1(n692), .Y(n82) );
  OAI22X1 U550 ( .A0(b[0]), .A1(n683), .B0(n693), .B1(n685), .Y(n395) );
  OAI22X1 U551 ( .A0(n693), .A1(n683), .B0(n694), .B1(n685), .Y(n394) );
  XNOR2X1 U552 ( .A(b[1]), .B(n647), .Y(n693) );
  OAI22X1 U553 ( .A0(n694), .A1(n683), .B0(n695), .B1(n685), .Y(n393) );
  XNOR2X1 U554 ( .A(b[2]), .B(n647), .Y(n694) );
  OAI22X1 U555 ( .A0(n695), .A1(n683), .B0(n696), .B1(n685), .Y(n392) );
  XNOR2X1 U556 ( .A(b[3]), .B(n647), .Y(n695) );
  OAI22X1 U557 ( .A0(n696), .A1(n683), .B0(n697), .B1(n685), .Y(n391) );
  XNOR2X1 U558 ( .A(b[4]), .B(n647), .Y(n696) );
  OAI22X1 U559 ( .A0(n697), .A1(n683), .B0(n698), .B1(n685), .Y(n390) );
  XNOR2X1 U560 ( .A(b[5]), .B(n647), .Y(n697) );
  OAI22X1 U561 ( .A0(n698), .A1(n683), .B0(n699), .B1(n685), .Y(n389) );
  XNOR2X1 U562 ( .A(b[6]), .B(n647), .Y(n698) );
  OAI22X1 U563 ( .A0(n699), .A1(n683), .B0(n700), .B1(n685), .Y(n388) );
  XNOR2X1 U564 ( .A(b[7]), .B(n647), .Y(n699) );
  OAI22X1 U565 ( .A0(n700), .A1(n683), .B0(n701), .B1(n685), .Y(n387) );
  XNOR2X1 U566 ( .A(b[8]), .B(n647), .Y(n700) );
  OAI22X1 U567 ( .A0(n701), .A1(n683), .B0(n702), .B1(n685), .Y(n386) );
  XNOR2X1 U568 ( .A(b[9]), .B(n647), .Y(n701) );
  OAI22X1 U569 ( .A0(n702), .A1(n683), .B0(n703), .B1(n685), .Y(n385) );
  XNOR2X1 U570 ( .A(b[10]), .B(n647), .Y(n702) );
  OAI22X1 U571 ( .A0(n703), .A1(n683), .B0(n704), .B1(n685), .Y(n384) );
  XNOR2X1 U572 ( .A(b[11]), .B(n647), .Y(n703) );
  OAI22X1 U573 ( .A0(n704), .A1(n683), .B0(n705), .B1(n685), .Y(n383) );
  XNOR2X1 U574 ( .A(b[12]), .B(n647), .Y(n704) );
  OAI22X1 U575 ( .A0(n705), .A1(n683), .B0(n706), .B1(n685), .Y(n382) );
  XNOR2X1 U576 ( .A(b[13]), .B(n647), .Y(n705) );
  OAI2BB2X1 U577 ( .B0(n706), .B1(n683), .A0N(n707), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U578 ( .A(b[14]), .B(n647), .Y(n706) );
  AOI22X1 U579 ( .A0(a[0]), .A1(n707), .B0(n708), .B1(n707), .Y(n380) );
  XNOR2X1 U580 ( .A(b[15]), .B(n684), .Y(n707) );
  NOR2X1 U581 ( .A(n709), .B(n686), .Y(n379) );
  OAI22X1 U582 ( .A0(n710), .A1(n711), .B0(n709), .B1(n712), .Y(n378) );
  XNOR2X1 U583 ( .A(n648), .B(b[0]), .Y(n710) );
  OAI22X1 U584 ( .A0(n712), .A1(n711), .B0(n709), .B1(n713), .Y(n377) );
  XNOR2X1 U585 ( .A(b[1]), .B(n648), .Y(n712) );
  OAI22X1 U586 ( .A0(n713), .A1(n711), .B0(n709), .B1(n714), .Y(n376) );
  XNOR2X1 U587 ( .A(b[2]), .B(n648), .Y(n713) );
  OAI22X1 U588 ( .A0(n714), .A1(n711), .B0(n709), .B1(n715), .Y(n375) );
  XNOR2X1 U589 ( .A(b[3]), .B(n648), .Y(n714) );
  OAI22X1 U590 ( .A0(n715), .A1(n711), .B0(n709), .B1(n716), .Y(n374) );
  XNOR2X1 U591 ( .A(b[4]), .B(n648), .Y(n715) );
  OAI22X1 U592 ( .A0(n716), .A1(n711), .B0(n709), .B1(n717), .Y(n373) );
  XNOR2X1 U593 ( .A(b[5]), .B(n648), .Y(n716) );
  OAI22X1 U594 ( .A0(n717), .A1(n711), .B0(n709), .B1(n718), .Y(n372) );
  XNOR2X1 U595 ( .A(b[6]), .B(n648), .Y(n717) );
  OAI22X1 U596 ( .A0(n718), .A1(n711), .B0(n709), .B1(n719), .Y(n371) );
  XNOR2X1 U597 ( .A(b[7]), .B(n648), .Y(n718) );
  OAI22X1 U598 ( .A0(n719), .A1(n711), .B0(n709), .B1(n720), .Y(n370) );
  XNOR2X1 U599 ( .A(b[8]), .B(n648), .Y(n719) );
  OAI22X1 U600 ( .A0(n720), .A1(n711), .B0(n709), .B1(n721), .Y(n369) );
  XNOR2X1 U601 ( .A(b[9]), .B(n648), .Y(n720) );
  OAI22X1 U602 ( .A0(n721), .A1(n711), .B0(n709), .B1(n722), .Y(n368) );
  XNOR2X1 U603 ( .A(b[10]), .B(n648), .Y(n721) );
  OAI22X1 U604 ( .A0(n722), .A1(n711), .B0(n709), .B1(n723), .Y(n367) );
  XNOR2X1 U605 ( .A(b[11]), .B(n648), .Y(n722) );
  OAI22X1 U606 ( .A0(n723), .A1(n711), .B0(n709), .B1(n724), .Y(n366) );
  XNOR2X1 U607 ( .A(b[12]), .B(n648), .Y(n723) );
  OAI2BB2X1 U608 ( .B0(n724), .B1(n711), .A0N(n682), .A1N(n725), .Y(n365) );
  XNOR2X1 U609 ( .A(b[13]), .B(n648), .Y(n724) );
  AOI22X1 U610 ( .A0(n726), .A1(n682), .B0(n680), .B1(n726), .Y(n364) );
  NOR2X1 U611 ( .A(n727), .B(n686), .Y(n363) );
  OAI22X1 U612 ( .A0(n728), .A1(n729), .B0(n727), .B1(n730), .Y(n362) );
  XNOR2X1 U613 ( .A(n649), .B(b[0]), .Y(n728) );
  OAI22X1 U614 ( .A0(n730), .A1(n729), .B0(n727), .B1(n731), .Y(n361) );
  XNOR2X1 U615 ( .A(b[1]), .B(n649), .Y(n730) );
  OAI22X1 U616 ( .A0(n731), .A1(n729), .B0(n727), .B1(n732), .Y(n360) );
  XNOR2X1 U617 ( .A(b[2]), .B(n649), .Y(n731) );
  OAI22X1 U618 ( .A0(n732), .A1(n729), .B0(n727), .B1(n733), .Y(n359) );
  XNOR2X1 U619 ( .A(b[3]), .B(n649), .Y(n732) );
  OAI22X1 U620 ( .A0(n733), .A1(n729), .B0(n727), .B1(n734), .Y(n358) );
  XNOR2X1 U621 ( .A(b[4]), .B(n649), .Y(n733) );
  OAI22X1 U622 ( .A0(n734), .A1(n729), .B0(n727), .B1(n735), .Y(n357) );
  XNOR2X1 U623 ( .A(b[5]), .B(n649), .Y(n734) );
  OAI22X1 U624 ( .A0(n735), .A1(n729), .B0(n727), .B1(n736), .Y(n356) );
  XNOR2X1 U625 ( .A(b[6]), .B(n649), .Y(n735) );
  OAI22X1 U626 ( .A0(n736), .A1(n729), .B0(n727), .B1(n737), .Y(n355) );
  XNOR2X1 U627 ( .A(b[7]), .B(n649), .Y(n736) );
  OAI22X1 U628 ( .A0(n737), .A1(n729), .B0(n727), .B1(n738), .Y(n354) );
  XNOR2X1 U629 ( .A(b[8]), .B(n649), .Y(n737) );
  OAI22X1 U630 ( .A0(n738), .A1(n729), .B0(n727), .B1(n739), .Y(n353) );
  XNOR2X1 U631 ( .A(b[9]), .B(n649), .Y(n738) );
  OAI22X1 U632 ( .A0(n739), .A1(n729), .B0(n727), .B1(n740), .Y(n352) );
  XNOR2X1 U633 ( .A(b[10]), .B(n649), .Y(n739) );
  OAI22X1 U634 ( .A0(n740), .A1(n729), .B0(n727), .B1(n741), .Y(n351) );
  XNOR2X1 U635 ( .A(b[11]), .B(n649), .Y(n740) );
  OAI22X1 U636 ( .A0(n741), .A1(n729), .B0(n727), .B1(n742), .Y(n350) );
  XNOR2X1 U637 ( .A(b[12]), .B(n649), .Y(n741) );
  OAI2BB2X1 U638 ( .B0(n742), .B1(n729), .A0N(n678), .A1N(n743), .Y(n349) );
  XNOR2X1 U639 ( .A(b[13]), .B(n649), .Y(n742) );
  AOI22X1 U640 ( .A0(n744), .A1(n678), .B0(n676), .B1(n744), .Y(n348) );
  NOR2X1 U641 ( .A(n745), .B(n686), .Y(n347) );
  OAI22X1 U642 ( .A0(n746), .A1(n747), .B0(n745), .B1(n748), .Y(n346) );
  XNOR2X1 U643 ( .A(n650), .B(b[0]), .Y(n746) );
  OAI22X1 U644 ( .A0(n748), .A1(n747), .B0(n745), .B1(n749), .Y(n345) );
  XNOR2X1 U645 ( .A(b[1]), .B(n650), .Y(n748) );
  OAI22X1 U646 ( .A0(n749), .A1(n747), .B0(n745), .B1(n750), .Y(n344) );
  XNOR2X1 U647 ( .A(b[2]), .B(n650), .Y(n749) );
  OAI22X1 U648 ( .A0(n750), .A1(n747), .B0(n745), .B1(n751), .Y(n343) );
  XNOR2X1 U649 ( .A(b[3]), .B(n650), .Y(n750) );
  OAI22X1 U650 ( .A0(n751), .A1(n747), .B0(n745), .B1(n752), .Y(n342) );
  XNOR2X1 U651 ( .A(b[4]), .B(n650), .Y(n751) );
  OAI22X1 U652 ( .A0(n752), .A1(n747), .B0(n745), .B1(n753), .Y(n341) );
  XNOR2X1 U653 ( .A(b[5]), .B(n650), .Y(n752) );
  OAI22X1 U654 ( .A0(n753), .A1(n747), .B0(n745), .B1(n754), .Y(n340) );
  XNOR2X1 U655 ( .A(b[6]), .B(n650), .Y(n753) );
  OAI22X1 U656 ( .A0(n754), .A1(n747), .B0(n745), .B1(n755), .Y(n339) );
  XNOR2X1 U657 ( .A(b[7]), .B(n650), .Y(n754) );
  OAI22X1 U658 ( .A0(n755), .A1(n747), .B0(n745), .B1(n756), .Y(n338) );
  XNOR2X1 U659 ( .A(b[8]), .B(n650), .Y(n755) );
  OAI22X1 U660 ( .A0(n757), .A1(n747), .B0(n745), .B1(n758), .Y(n336) );
  OAI22X1 U661 ( .A0(n758), .A1(n747), .B0(n745), .B1(n759), .Y(n335) );
  XNOR2X1 U662 ( .A(b[11]), .B(n650), .Y(n758) );
  OAI22X1 U663 ( .A0(n759), .A1(n747), .B0(n745), .B1(n760), .Y(n334) );
  XNOR2X1 U664 ( .A(b[12]), .B(n650), .Y(n759) );
  OAI22X1 U665 ( .A0(n760), .A1(n747), .B0(n745), .B1(n761), .Y(n333) );
  XNOR2X1 U666 ( .A(b[13]), .B(n650), .Y(n760) );
  OAI2BB2X1 U667 ( .B0(n761), .B1(n747), .A0N(n674), .A1N(n762), .Y(n332) );
  XNOR2X1 U668 ( .A(b[14]), .B(n650), .Y(n761) );
  AOI22X1 U669 ( .A0(n762), .A1(n674), .B0(n672), .B1(n762), .Y(n331) );
  XNOR2X1 U670 ( .A(b[15]), .B(n673), .Y(n762) );
  NOR2X1 U671 ( .A(n763), .B(n686), .Y(n330) );
  OAI22X1 U672 ( .A0(n764), .A1(n765), .B0(n763), .B1(n766), .Y(n329) );
  XNOR2X1 U673 ( .A(n651), .B(b[0]), .Y(n764) );
  OAI22X1 U674 ( .A0(n766), .A1(n765), .B0(n763), .B1(n767), .Y(n328) );
  XNOR2X1 U675 ( .A(b[1]), .B(n651), .Y(n766) );
  OAI22X1 U676 ( .A0(n767), .A1(n765), .B0(n763), .B1(n768), .Y(n327) );
  XNOR2X1 U677 ( .A(b[2]), .B(n651), .Y(n767) );
  OAI22X1 U678 ( .A0(n768), .A1(n765), .B0(n763), .B1(n769), .Y(n326) );
  XNOR2X1 U679 ( .A(b[3]), .B(n651), .Y(n768) );
  OAI22X1 U680 ( .A0(n769), .A1(n765), .B0(n763), .B1(n770), .Y(n325) );
  XNOR2X1 U681 ( .A(b[4]), .B(n651), .Y(n769) );
  OAI22X1 U682 ( .A0(n770), .A1(n765), .B0(n763), .B1(n771), .Y(n324) );
  XNOR2X1 U683 ( .A(b[5]), .B(n651), .Y(n770) );
  OAI22X1 U684 ( .A0(n771), .A1(n765), .B0(n763), .B1(n772), .Y(n323) );
  XNOR2X1 U685 ( .A(b[6]), .B(n651), .Y(n771) );
  OAI22X1 U686 ( .A0(n772), .A1(n765), .B0(n763), .B1(n773), .Y(n322) );
  XNOR2X1 U687 ( .A(b[7]), .B(n651), .Y(n772) );
  OAI22X1 U688 ( .A0(n773), .A1(n765), .B0(n763), .B1(n774), .Y(n321) );
  XNOR2X1 U689 ( .A(b[8]), .B(n651), .Y(n773) );
  OAI22X1 U690 ( .A0(n774), .A1(n765), .B0(n763), .B1(n775), .Y(n320) );
  XNOR2X1 U691 ( .A(b[9]), .B(n651), .Y(n774) );
  OAI22X1 U692 ( .A0(n775), .A1(n765), .B0(n763), .B1(n776), .Y(n319) );
  XNOR2X1 U693 ( .A(b[10]), .B(n651), .Y(n775) );
  OAI22X1 U694 ( .A0(n776), .A1(n765), .B0(n763), .B1(n777), .Y(n318) );
  XNOR2X1 U695 ( .A(b[11]), .B(n651), .Y(n776) );
  OAI22X1 U696 ( .A0(n777), .A1(n765), .B0(n763), .B1(n778), .Y(n317) );
  XNOR2X1 U697 ( .A(b[12]), .B(n651), .Y(n777) );
  OAI2BB2X1 U698 ( .B0(n778), .B1(n765), .A0N(n671), .A1N(n779), .Y(n316) );
  XNOR2X1 U699 ( .A(b[13]), .B(n651), .Y(n778) );
  AOI22X1 U700 ( .A0(n780), .A1(n671), .B0(n669), .B1(n780), .Y(n315) );
  NOR2X1 U701 ( .A(n781), .B(n686), .Y(n314) );
  OAI22X1 U702 ( .A0(n782), .A1(n783), .B0(n781), .B1(n784), .Y(n313) );
  XNOR2X1 U703 ( .A(n652), .B(b[0]), .Y(n782) );
  OAI22X1 U704 ( .A0(n784), .A1(n783), .B0(n781), .B1(n785), .Y(n312) );
  XNOR2X1 U705 ( .A(b[1]), .B(n652), .Y(n784) );
  OAI22X1 U706 ( .A0(n785), .A1(n783), .B0(n781), .B1(n786), .Y(n311) );
  XNOR2X1 U707 ( .A(b[2]), .B(n652), .Y(n785) );
  OAI22X1 U708 ( .A0(n786), .A1(n783), .B0(n781), .B1(n787), .Y(n310) );
  XNOR2X1 U709 ( .A(b[3]), .B(n652), .Y(n786) );
  OAI22X1 U710 ( .A0(n787), .A1(n783), .B0(n781), .B1(n788), .Y(n309) );
  XNOR2X1 U711 ( .A(b[4]), .B(n652), .Y(n787) );
  OAI22X1 U712 ( .A0(n788), .A1(n783), .B0(n781), .B1(n789), .Y(n308) );
  XNOR2X1 U713 ( .A(b[5]), .B(n652), .Y(n788) );
  OAI22X1 U714 ( .A0(n789), .A1(n783), .B0(n781), .B1(n790), .Y(n307) );
  XNOR2X1 U715 ( .A(b[6]), .B(n652), .Y(n789) );
  OAI22X1 U716 ( .A0(n790), .A1(n783), .B0(n781), .B1(n791), .Y(n306) );
  XNOR2X1 U717 ( .A(b[7]), .B(n652), .Y(n790) );
  OAI22X1 U718 ( .A0(n791), .A1(n783), .B0(n781), .B1(n792), .Y(n305) );
  XNOR2X1 U719 ( .A(b[8]), .B(n652), .Y(n791) );
  OAI22X1 U720 ( .A0(n792), .A1(n783), .B0(n781), .B1(n793), .Y(n304) );
  XNOR2X1 U721 ( .A(b[9]), .B(n652), .Y(n792) );
  OAI22X1 U722 ( .A0(n794), .A1(n783), .B0(n781), .B1(n795), .Y(n303) );
  OAI22X1 U723 ( .A0(n795), .A1(n783), .B0(n781), .B1(n796), .Y(n302) );
  XNOR2X1 U724 ( .A(b[12]), .B(n652), .Y(n795) );
  OAI2BB2X1 U725 ( .B0(n796), .B1(n783), .A0N(n667), .A1N(n687), .Y(n301) );
  XOR2X1 U726 ( .A(b[14]), .B(n652), .Y(n687) );
  XNOR2X1 U727 ( .A(b[13]), .B(n652), .Y(n796) );
  AOI22X1 U728 ( .A0(n688), .A1(n667), .B0(n665), .B1(n688), .Y(n300) );
  XNOR2X1 U729 ( .A(b[15]), .B(n666), .Y(n688) );
  NOR2X1 U730 ( .A(n797), .B(n686), .Y(n299) );
  OAI22X1 U731 ( .A0(n798), .A1(n799), .B0(n797), .B1(n800), .Y(n298) );
  XNOR2X1 U732 ( .A(n653), .B(b[0]), .Y(n798) );
  OAI22X1 U733 ( .A0(n800), .A1(n799), .B0(n797), .B1(n801), .Y(n297) );
  XNOR2X1 U734 ( .A(b[1]), .B(n653), .Y(n800) );
  OAI22X1 U735 ( .A0(n801), .A1(n799), .B0(n797), .B1(n802), .Y(n296) );
  XNOR2X1 U736 ( .A(b[2]), .B(n653), .Y(n801) );
  OAI22X1 U737 ( .A0(n803), .A1(n799), .B0(n797), .B1(n804), .Y(n294) );
  OAI22X1 U738 ( .A0(n804), .A1(n799), .B0(n797), .B1(n805), .Y(n293) );
  XNOR2X1 U739 ( .A(b[5]), .B(n653), .Y(n804) );
  OAI22X1 U740 ( .A0(n805), .A1(n799), .B0(n797), .B1(n806), .Y(n292) );
  XNOR2X1 U741 ( .A(b[6]), .B(n653), .Y(n805) );
  OAI22X1 U742 ( .A0(n806), .A1(n799), .B0(n797), .B1(n807), .Y(n291) );
  XNOR2X1 U743 ( .A(b[7]), .B(n653), .Y(n806) );
  OAI22X1 U744 ( .A0(n807), .A1(n799), .B0(n797), .B1(n808), .Y(n290) );
  XNOR2X1 U745 ( .A(b[8]), .B(n653), .Y(n807) );
  OAI22X1 U746 ( .A0(n808), .A1(n799), .B0(n797), .B1(n809), .Y(n289) );
  XNOR2X1 U747 ( .A(b[9]), .B(n653), .Y(n808) );
  OAI22X1 U748 ( .A0(n809), .A1(n799), .B0(n797), .B1(n810), .Y(n288) );
  XNOR2X1 U749 ( .A(b[10]), .B(n653), .Y(n809) );
  OAI22X1 U750 ( .A0(n810), .A1(n799), .B0(n797), .B1(n811), .Y(n287) );
  XNOR2X1 U751 ( .A(b[11]), .B(n653), .Y(n810) );
  OAI22X1 U752 ( .A0(n811), .A1(n799), .B0(n797), .B1(n812), .Y(n286) );
  XNOR2X1 U753 ( .A(b[12]), .B(n653), .Y(n811) );
  OAI2BB2X1 U754 ( .B0(n812), .B1(n799), .A0N(n662), .A1N(n689), .Y(n285) );
  XOR2X1 U755 ( .A(b[14]), .B(n653), .Y(n689) );
  XNOR2X1 U756 ( .A(b[13]), .B(n653), .Y(n812) );
  AOI22X1 U757 ( .A0(n690), .A1(n662), .B0(n660), .B1(n690), .Y(n284) );
  XNOR2X1 U758 ( .A(b[15]), .B(n661), .Y(n690) );
  NOR2X1 U759 ( .A(n813), .B(n686), .Y(n283) );
  OAI22X1 U760 ( .A0(n814), .A1(n815), .B0(n813), .B1(n816), .Y(n282) );
  XNOR2X1 U761 ( .A(n654), .B(b[0]), .Y(n814) );
  OAI22X1 U762 ( .A0(n816), .A1(n815), .B0(n813), .B1(n817), .Y(n281) );
  XNOR2X1 U763 ( .A(b[1]), .B(n654), .Y(n816) );
  OAI22X1 U764 ( .A0(n817), .A1(n815), .B0(n813), .B1(n818), .Y(n280) );
  XNOR2X1 U765 ( .A(b[2]), .B(n654), .Y(n817) );
  OAI22X1 U766 ( .A0(n818), .A1(n815), .B0(n813), .B1(n819), .Y(n279) );
  XNOR2X1 U767 ( .A(b[3]), .B(n654), .Y(n818) );
  OAI22X1 U768 ( .A0(n819), .A1(n815), .B0(n813), .B1(n820), .Y(n278) );
  XNOR2X1 U769 ( .A(b[4]), .B(n654), .Y(n819) );
  OAI22X1 U770 ( .A0(n820), .A1(n815), .B0(n813), .B1(n821), .Y(n277) );
  XNOR2X1 U771 ( .A(b[5]), .B(n654), .Y(n820) );
  OAI22X1 U772 ( .A0(n821), .A1(n815), .B0(n813), .B1(n822), .Y(n276) );
  XNOR2X1 U773 ( .A(b[6]), .B(n654), .Y(n821) );
  OAI22X1 U774 ( .A0(n822), .A1(n815), .B0(n813), .B1(n823), .Y(n275) );
  XNOR2X1 U775 ( .A(b[7]), .B(n654), .Y(n822) );
  OAI22X1 U776 ( .A0(n823), .A1(n815), .B0(n813), .B1(n824), .Y(n274) );
  XNOR2X1 U777 ( .A(b[8]), .B(n654), .Y(n823) );
  OAI22X1 U778 ( .A0(n824), .A1(n815), .B0(n813), .B1(n825), .Y(n273) );
  XNOR2X1 U779 ( .A(b[9]), .B(n654), .Y(n824) );
  OAI22X1 U780 ( .A0(n825), .A1(n815), .B0(n813), .B1(n826), .Y(n272) );
  XNOR2X1 U781 ( .A(b[10]), .B(n654), .Y(n825) );
  OAI22X1 U782 ( .A0(n826), .A1(n815), .B0(n813), .B1(n827), .Y(n271) );
  XNOR2X1 U783 ( .A(b[11]), .B(n654), .Y(n826) );
  OAI22X1 U784 ( .A0(n827), .A1(n815), .B0(n813), .B1(n828), .Y(n270) );
  XNOR2X1 U785 ( .A(b[12]), .B(n654), .Y(n827) );
  OAI2BB2X1 U786 ( .B0(n828), .B1(n815), .A0N(n658), .A1N(n691), .Y(n269) );
  XOR2X1 U787 ( .A(b[14]), .B(n654), .Y(n691) );
  XNOR2X1 U788 ( .A(b[13]), .B(n654), .Y(n828) );
  AOI22X1 U789 ( .A0(n692), .A1(n658), .B0(n656), .B1(n692), .Y(n268) );
  XNOR2X1 U790 ( .A(b[15]), .B(n657), .Y(n692) );
  OAI21XL U791 ( .A0(b[0]), .A1(n684), .B0(n683), .Y(n267) );
  NOR2X1 U792 ( .A(n684), .B(a[0]), .Y(n708) );
  OAI32X1 U793 ( .A0(n681), .A1(b[0]), .A2(n709), .B0(n681), .B1(n711), .Y(
        n266) );
  OAI32X1 U794 ( .A0(n677), .A1(b[0]), .A2(n727), .B0(n677), .B1(n729), .Y(
        n265) );
  OAI32X1 U795 ( .A0(n673), .A1(b[0]), .A2(n745), .B0(n673), .B1(n747), .Y(
        n264) );
  OAI32X1 U796 ( .A0(n670), .A1(b[0]), .A2(n763), .B0(n670), .B1(n765), .Y(
        n263) );
  OAI32X1 U797 ( .A0(n666), .A1(b[0]), .A2(n781), .B0(n666), .B1(n783), .Y(
        n262) );
  OAI32X1 U798 ( .A0(n661), .A1(b[0]), .A2(n797), .B0(n661), .B1(n799), .Y(
        n261) );
  OAI32X1 U799 ( .A0(n657), .A1(b[0]), .A2(n813), .B0(n657), .B1(n815), .Y(
        n260) );
  XNOR2X1 U800 ( .A(n657), .B(a[14]), .Y(n829) );
  XNOR2X1 U801 ( .A(n830), .B(n831), .Y(n171) );
  OR2X1 U802 ( .A(n830), .B(n831), .Y(n170) );
  OAI22X1 U803 ( .A0(n756), .A1(n747), .B0(n745), .B1(n757), .Y(n831) );
  XNOR2X1 U804 ( .A(b[10]), .B(n650), .Y(n757) );
  XNOR2X1 U805 ( .A(n673), .B(a[6]), .Y(n832) );
  XNOR2X1 U806 ( .A(b[9]), .B(n650), .Y(n756) );
  OAI22X1 U807 ( .A0(n802), .A1(n799), .B0(n797), .B1(n803), .Y(n830) );
  XNOR2X1 U808 ( .A(b[4]), .B(n653), .Y(n803) );
  XNOR2X1 U809 ( .A(n661), .B(a[12]), .Y(n833) );
  XNOR2X1 U810 ( .A(b[3]), .B(n653), .Y(n802) );
  AOI22X1 U811 ( .A0(n725), .A1(n680), .B0(n682), .B1(n726), .Y(n160) );
  XNOR2X1 U812 ( .A(b[15]), .B(n681), .Y(n726) );
  XNOR2X1 U813 ( .A(n681), .B(a[2]), .Y(n834) );
  XOR2X1 U814 ( .A(b[14]), .B(n648), .Y(n725) );
  AOI22X1 U815 ( .A0(n743), .A1(n676), .B0(n678), .B1(n744), .Y(n140) );
  XNOR2X1 U816 ( .A(b[15]), .B(n677), .Y(n744) );
  XNOR2X1 U817 ( .A(n677), .B(a[4]), .Y(n835) );
  XOR2X1 U818 ( .A(b[14]), .B(n649), .Y(n743) );
  OAI22X1 U819 ( .A0(n793), .A1(n783), .B0(n781), .B1(n794), .Y(n121) );
  XNOR2X1 U820 ( .A(b[11]), .B(n652), .Y(n794) );
  XNOR2X1 U821 ( .A(n666), .B(a[10]), .Y(n836) );
  XNOR2X1 U822 ( .A(b[10]), .B(n652), .Y(n793) );
  AOI22X1 U823 ( .A0(n779), .A1(n669), .B0(n671), .B1(n780), .Y(n108) );
  XNOR2X1 U824 ( .A(b[15]), .B(n670), .Y(n780) );
  XNOR2X1 U825 ( .A(n670), .B(a[8]), .Y(n837) );
  XOR2X1 U826 ( .A(b[14]), .B(n651), .Y(n779) );
endmodule


module PE_56 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_56_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_56_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_56_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_56_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n658), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n657), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n656), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n661), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n662), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n660), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n659), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n659) );
  INVX1 U492 ( .A(n121), .Y(n662) );
  INVX1 U493 ( .A(n96), .Y(n656) );
  INVX1 U494 ( .A(n82), .Y(n658) );
  INVX1 U495 ( .A(n648), .Y(n679) );
  CLKINVX3 U496 ( .A(n709), .Y(n678) );
  CLKINVX3 U497 ( .A(n651), .Y(n670) );
  CLKINVX3 U498 ( .A(n649), .Y(n676) );
  CLKINVX3 U499 ( .A(n650), .Y(n673) );
  CLKINVX3 U500 ( .A(n647), .Y(n663) );
  CLKINVX3 U501 ( .A(n652), .Y(n667) );
  CLKINVX3 U502 ( .A(n653), .Y(n686) );
  CLKINVX3 U503 ( .A(n654), .Y(n684) );
  INVX1 U504 ( .A(n655), .Y(n681) );
  INVX1 U505 ( .A(n728), .Y(n674) );
  INVX1 U506 ( .A(n710), .Y(n677) );
  INVX1 U507 ( .A(n712), .Y(n675) );
  INVX1 U508 ( .A(n730), .Y(n672) );
  INVX1 U509 ( .A(n140), .Y(n660) );
  INVX1 U510 ( .A(n764), .Y(n668) );
  INVX1 U511 ( .A(n746), .Y(n671) );
  INVX1 U512 ( .A(n748), .Y(n669) );
  INVX1 U513 ( .A(n108), .Y(n661) );
  INVX1 U514 ( .A(n782), .Y(n666) );
  INVX1 U515 ( .A(n766), .Y(n664) );
  INVX1 U516 ( .A(n784), .Y(n665) );
  INVX1 U517 ( .A(n798), .Y(n685) );
  INVX1 U518 ( .A(n88), .Y(n657) );
  INVX1 U519 ( .A(n814), .Y(n682) );
  INVX1 U520 ( .A(n800), .Y(n683) );
  INVX1 U521 ( .A(n816), .Y(n680) );
  XOR2X2 U522 ( .A(a[2]), .B(n679), .Y(n710) );
  BUFX3 U523 ( .A(a[1]), .Y(n648) );
  XOR2X2 U524 ( .A(a[6]), .B(n673), .Y(n746) );
  XOR2X2 U525 ( .A(a[4]), .B(n676), .Y(n728) );
  XOR2X2 U526 ( .A(a[8]), .B(n670), .Y(n764) );
  CLKINVX3 U527 ( .A(a[0]), .Y(n687) );
  BUFX3 U528 ( .A(b[0]), .Y(n647) );
  BUFX3 U529 ( .A(a[7]), .Y(n651) );
  BUFX3 U530 ( .A(a[3]), .Y(n649) );
  BUFX3 U531 ( .A(a[5]), .Y(n650) );
  XOR2X2 U532 ( .A(a[10]), .B(n667), .Y(n782) );
  XOR2X2 U533 ( .A(a[12]), .B(n686), .Y(n798) );
  BUFX3 U534 ( .A(a[9]), .Y(n652) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n684), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n687), .B(n663), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n665), .B0(n666), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n683), .B0(n685), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n680), .B0(n682), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n678), .B0(n694), .B1(n687), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n678), .B0(n695), .B1(n687), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n678), .B0(n696), .B1(n687), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n678), .B0(n697), .B1(n687), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n678), .B0(n698), .B1(n687), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n678), .B0(n699), .B1(n687), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n678), .B0(n700), .B1(n687), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n678), .B0(n701), .B1(n687), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n678), .B0(n702), .B1(n687), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n678), .B0(n703), .B1(n687), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n678), .B0(n704), .B1(n687), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n678), .B0(n705), .B1(n687), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n678), .B0(n706), .B1(n687), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n678), .B0(n707), .B1(n687), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n678), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n679), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n663), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n677), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n677), .B0(n675), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n663), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n674), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n674), .B0(n672), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n663), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n671), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n671), .B0(n669), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n670), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n663), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n668), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n668), .B0(n664), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n663), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n666), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n666), .B0(n665), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n686), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n663), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n685), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n685), .B0(n683), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n684), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n663), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n682), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n682), .B0(n680), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n681), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n679), .B0(n678), .Y(n267) );
  NOR2X1 U793 ( .A(n679), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n676), .A1(n647), .A2(n710), .B0(n676), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n673), .A1(n647), .A2(n728), .B0(n673), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n670), .A1(n647), .A2(n746), .B0(n670), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n667), .A1(n647), .A2(n764), .B0(n667), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n686), .A1(n647), .A2(n782), .B0(n686), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n684), .A1(n647), .A2(n798), .B0(n684), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n681), .A1(n647), .A2(n814), .B0(n681), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n681), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n670), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n684), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n675), .B0(n677), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n676), .Y(n727) );
  XNOR2X1 U814 ( .A(n676), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n672), .B0(n674), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n673), .Y(n745) );
  XNOR2X1 U818 ( .A(n673), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n686), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n664), .B0(n668), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n667), .Y(n781) );
  XNOR2X1 U826 ( .A(n667), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_57 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_57_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_57_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_57_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_57_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  CLKINVX3 U495 ( .A(n709), .Y(n684) );
  CLKINVX3 U496 ( .A(n649), .Y(n682) );
  INVX1 U497 ( .A(n648), .Y(n685) );
  CLKINVX3 U498 ( .A(n651), .Y(n674) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n652), .Y(n671) );
  CLKINVX3 U501 ( .A(n647), .Y(n687) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n710), .Y(n683) );
  INVX1 U505 ( .A(n712), .Y(n681) );
  INVX1 U506 ( .A(n655), .Y(n658) );
  INVX1 U507 ( .A(n728), .Y(n679) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n746), .Y(n675) );
  INVX1 U511 ( .A(n764), .Y(n672) );
  INVX1 U512 ( .A(n766), .Y(n670) );
  INVX1 U513 ( .A(n748), .Y(n673) );
  INVX1 U514 ( .A(n108), .Y(n669) );
  INVX1 U515 ( .A(n782), .Y(n668) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n800), .Y(n661) );
  INVX1 U519 ( .A(n88), .Y(n660) );
  INVX1 U520 ( .A(n814), .Y(n659) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U523 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U524 ( .A(a[3]), .Y(n649) );
  BUFX3 U525 ( .A(a[1]), .Y(n648) );
  XOR2X2 U526 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U527 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U528 ( .A(a[0]), .Y(n686) );
  BUFX3 U529 ( .A(a[7]), .Y(n651) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(a[9]), .Y(n652) );
  BUFX3 U532 ( .A(b[0]), .Y(n647) );
  XOR2X2 U533 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U534 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_58 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_58_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_58_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_58_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_58_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  CLKINVX3 U495 ( .A(n709), .Y(n684) );
  CLKINVX3 U496 ( .A(n649), .Y(n682) );
  INVX1 U497 ( .A(n648), .Y(n685) );
  CLKINVX3 U498 ( .A(n651), .Y(n674) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n652), .Y(n671) );
  CLKINVX3 U501 ( .A(n647), .Y(n687) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n710), .Y(n683) );
  INVX1 U505 ( .A(n712), .Y(n681) );
  INVX1 U506 ( .A(n655), .Y(n658) );
  INVX1 U507 ( .A(n728), .Y(n679) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n746), .Y(n675) );
  INVX1 U511 ( .A(n764), .Y(n672) );
  INVX1 U512 ( .A(n766), .Y(n670) );
  INVX1 U513 ( .A(n748), .Y(n673) );
  INVX1 U514 ( .A(n108), .Y(n669) );
  INVX1 U515 ( .A(n782), .Y(n668) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n800), .Y(n661) );
  INVX1 U519 ( .A(n88), .Y(n660) );
  INVX1 U520 ( .A(n814), .Y(n659) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U523 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U524 ( .A(a[3]), .Y(n649) );
  BUFX3 U525 ( .A(a[1]), .Y(n648) );
  XOR2X2 U526 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U527 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U528 ( .A(a[0]), .Y(n686) );
  BUFX3 U529 ( .A(a[7]), .Y(n651) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(a[9]), .Y(n652) );
  BUFX3 U532 ( .A(b[0]), .Y(n647) );
  XOR2X2 U533 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U534 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_59 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_59_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_59_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_59_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_59_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  CLKINVX3 U495 ( .A(n709), .Y(n684) );
  CLKINVX3 U496 ( .A(n649), .Y(n682) );
  INVX1 U497 ( .A(n648), .Y(n685) );
  CLKINVX3 U498 ( .A(n651), .Y(n674) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n652), .Y(n671) );
  CLKINVX3 U501 ( .A(n647), .Y(n687) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n710), .Y(n683) );
  INVX1 U505 ( .A(n712), .Y(n681) );
  INVX1 U506 ( .A(n655), .Y(n658) );
  INVX1 U507 ( .A(n728), .Y(n679) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n746), .Y(n675) );
  INVX1 U511 ( .A(n764), .Y(n672) );
  INVX1 U512 ( .A(n766), .Y(n670) );
  INVX1 U513 ( .A(n748), .Y(n673) );
  INVX1 U514 ( .A(n108), .Y(n669) );
  INVX1 U515 ( .A(n782), .Y(n668) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n800), .Y(n661) );
  INVX1 U519 ( .A(n88), .Y(n660) );
  INVX1 U520 ( .A(n814), .Y(n659) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U523 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U524 ( .A(a[3]), .Y(n649) );
  BUFX3 U525 ( .A(a[1]), .Y(n648) );
  XOR2X2 U526 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U527 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U528 ( .A(a[0]), .Y(n686) );
  BUFX3 U529 ( .A(a[7]), .Y(n651) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(a[9]), .Y(n652) );
  BUFX3 U532 ( .A(b[0]), .Y(n647) );
  XOR2X2 U533 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U534 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_60 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_60_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_60_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_60_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_60_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  CLKINVX3 U495 ( .A(n709), .Y(n684) );
  CLKINVX3 U496 ( .A(n649), .Y(n682) );
  INVX1 U497 ( .A(n648), .Y(n685) );
  CLKINVX3 U498 ( .A(n651), .Y(n674) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n652), .Y(n671) );
  CLKINVX3 U501 ( .A(n647), .Y(n687) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n710), .Y(n683) );
  INVX1 U505 ( .A(n712), .Y(n681) );
  INVX1 U506 ( .A(n655), .Y(n658) );
  INVX1 U507 ( .A(n728), .Y(n679) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n746), .Y(n675) );
  INVX1 U511 ( .A(n764), .Y(n672) );
  INVX1 U512 ( .A(n766), .Y(n670) );
  INVX1 U513 ( .A(n748), .Y(n673) );
  INVX1 U514 ( .A(n108), .Y(n669) );
  INVX1 U515 ( .A(n782), .Y(n668) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n800), .Y(n661) );
  INVX1 U519 ( .A(n88), .Y(n660) );
  INVX1 U520 ( .A(n814), .Y(n659) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U523 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U524 ( .A(a[3]), .Y(n649) );
  BUFX3 U525 ( .A(a[1]), .Y(n648) );
  XOR2X2 U526 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U527 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U528 ( .A(a[0]), .Y(n686) );
  BUFX3 U529 ( .A(a[7]), .Y(n651) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(a[9]), .Y(n652) );
  BUFX3 U532 ( .A(b[0]), .Y(n647) );
  XOR2X2 U533 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U534 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_61 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_61_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_61_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_61_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_61_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  CLKINVX3 U495 ( .A(n709), .Y(n684) );
  CLKINVX3 U496 ( .A(n649), .Y(n682) );
  INVX1 U497 ( .A(n648), .Y(n685) );
  CLKINVX3 U498 ( .A(n651), .Y(n674) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n652), .Y(n671) );
  CLKINVX3 U501 ( .A(n647), .Y(n687) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n710), .Y(n683) );
  INVX1 U505 ( .A(n712), .Y(n681) );
  INVX1 U506 ( .A(n655), .Y(n658) );
  INVX1 U507 ( .A(n728), .Y(n679) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n746), .Y(n675) );
  INVX1 U511 ( .A(n764), .Y(n672) );
  INVX1 U512 ( .A(n766), .Y(n670) );
  INVX1 U513 ( .A(n748), .Y(n673) );
  INVX1 U514 ( .A(n108), .Y(n669) );
  INVX1 U515 ( .A(n782), .Y(n668) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n800), .Y(n661) );
  INVX1 U519 ( .A(n88), .Y(n660) );
  INVX1 U520 ( .A(n814), .Y(n659) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U523 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U524 ( .A(a[3]), .Y(n649) );
  BUFX3 U525 ( .A(a[1]), .Y(n648) );
  XOR2X2 U526 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U527 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U528 ( .A(a[0]), .Y(n686) );
  BUFX3 U529 ( .A(a[7]), .Y(n651) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(a[9]), .Y(n652) );
  BUFX3 U532 ( .A(b[0]), .Y(n647) );
  XOR2X2 U533 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U534 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_62 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_62_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_62_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_62_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_62_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  CLKINVX3 U495 ( .A(n709), .Y(n684) );
  CLKINVX3 U496 ( .A(n649), .Y(n682) );
  INVX1 U497 ( .A(n648), .Y(n685) );
  CLKINVX3 U498 ( .A(n651), .Y(n674) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n652), .Y(n671) );
  CLKINVX3 U501 ( .A(n647), .Y(n687) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n710), .Y(n683) );
  INVX1 U505 ( .A(n712), .Y(n681) );
  INVX1 U506 ( .A(n655), .Y(n658) );
  INVX1 U507 ( .A(n728), .Y(n679) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n746), .Y(n675) );
  INVX1 U511 ( .A(n764), .Y(n672) );
  INVX1 U512 ( .A(n766), .Y(n670) );
  INVX1 U513 ( .A(n748), .Y(n673) );
  INVX1 U514 ( .A(n108), .Y(n669) );
  INVX1 U515 ( .A(n782), .Y(n668) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n800), .Y(n661) );
  INVX1 U519 ( .A(n88), .Y(n660) );
  INVX1 U520 ( .A(n814), .Y(n659) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U523 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U524 ( .A(a[3]), .Y(n649) );
  BUFX3 U525 ( .A(a[1]), .Y(n648) );
  XOR2X2 U526 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U527 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U528 ( .A(a[0]), .Y(n686) );
  BUFX3 U529 ( .A(a[7]), .Y(n651) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(a[9]), .Y(n652) );
  BUFX3 U532 ( .A(b[0]), .Y(n647) );
  XOR2X2 U533 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U534 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_63 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_63_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_63_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_63_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_63_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n656), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n660), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n664), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n669), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n665), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n676), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n680), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n680) );
  INVX1 U492 ( .A(n121), .Y(n665) );
  INVX1 U493 ( .A(n96), .Y(n664) );
  INVX1 U494 ( .A(n82), .Y(n656) );
  CLKINVX3 U495 ( .A(n709), .Y(n684) );
  CLKINVX3 U496 ( .A(n649), .Y(n682) );
  INVX1 U497 ( .A(n648), .Y(n685) );
  CLKINVX3 U498 ( .A(n651), .Y(n674) );
  CLKINVX3 U499 ( .A(n650), .Y(n678) );
  CLKINVX3 U500 ( .A(n652), .Y(n671) );
  CLKINVX3 U501 ( .A(n647), .Y(n687) );
  CLKINVX3 U502 ( .A(n653), .Y(n667) );
  CLKINVX3 U503 ( .A(n654), .Y(n662) );
  INVX1 U504 ( .A(n710), .Y(n683) );
  INVX1 U505 ( .A(n712), .Y(n681) );
  INVX1 U506 ( .A(n655), .Y(n658) );
  INVX1 U507 ( .A(n728), .Y(n679) );
  INVX1 U508 ( .A(n730), .Y(n677) );
  INVX1 U509 ( .A(n140), .Y(n676) );
  INVX1 U510 ( .A(n746), .Y(n675) );
  INVX1 U511 ( .A(n764), .Y(n672) );
  INVX1 U512 ( .A(n766), .Y(n670) );
  INVX1 U513 ( .A(n748), .Y(n673) );
  INVX1 U514 ( .A(n108), .Y(n669) );
  INVX1 U515 ( .A(n782), .Y(n668) );
  INVX1 U516 ( .A(n784), .Y(n666) );
  INVX1 U517 ( .A(n798), .Y(n663) );
  INVX1 U518 ( .A(n800), .Y(n661) );
  INVX1 U519 ( .A(n88), .Y(n660) );
  INVX1 U520 ( .A(n814), .Y(n659) );
  INVX1 U521 ( .A(n816), .Y(n657) );
  XOR2X2 U522 ( .A(a[4]), .B(n682), .Y(n728) );
  XOR2X2 U523 ( .A(a[2]), .B(n685), .Y(n710) );
  BUFX3 U524 ( .A(a[3]), .Y(n649) );
  BUFX3 U525 ( .A(a[1]), .Y(n648) );
  XOR2X2 U526 ( .A(a[6]), .B(n678), .Y(n746) );
  XOR2X2 U527 ( .A(a[8]), .B(n674), .Y(n764) );
  CLKINVX3 U528 ( .A(a[0]), .Y(n686) );
  BUFX3 U529 ( .A(a[7]), .Y(n651) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(a[9]), .Y(n652) );
  BUFX3 U532 ( .A(b[0]), .Y(n647) );
  XOR2X2 U533 ( .A(a[10]), .B(n671), .Y(n782) );
  XOR2X2 U534 ( .A(a[12]), .B(n667), .Y(n798) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n662), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n686), .B(n687), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n666), .B0(n668), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n661), .B0(n663), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n657), .B0(n659), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n684), .B0(n694), .B1(n686), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n684), .B0(n695), .B1(n686), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n684), .B0(n696), .B1(n686), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n684), .B0(n697), .B1(n686), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n684), .B0(n698), .B1(n686), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n684), .B0(n699), .B1(n686), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n684), .B0(n700), .B1(n686), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n684), .B0(n701), .B1(n686), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n684), .B0(n702), .B1(n686), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n684), .B0(n703), .B1(n686), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n684), .B0(n704), .B1(n686), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n684), .B0(n705), .B1(n686), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n684), .B0(n706), .B1(n686), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n684), .B0(n707), .B1(n686), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n684), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n685), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n687), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n683), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n683), .B0(n681), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n687), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n679), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n679), .B0(n677), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n687), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n675), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n675), .B0(n673), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n674), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n687), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n672), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n672), .B0(n670), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n687), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n668), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n668), .B0(n666), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n667), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n687), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n663), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n663), .B0(n661), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n662), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n687), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n659), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n659), .B0(n657), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n658), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n685), .B0(n684), .Y(n267) );
  NOR2X1 U793 ( .A(n685), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n682), .A1(n647), .A2(n710), .B0(n682), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n678), .A1(n647), .A2(n728), .B0(n678), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n674), .A1(n647), .A2(n746), .B0(n674), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n671), .A1(n647), .A2(n764), .B0(n671), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n667), .A1(n647), .A2(n782), .B0(n667), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n662), .A1(n647), .A2(n798), .B0(n662), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n658), .A1(n647), .A2(n814), .B0(n658), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n658), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n674), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n662), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n681), .B0(n683), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n682), .Y(n727) );
  XNOR2X1 U814 ( .A(n682), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n677), .B0(n679), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n678), .Y(n745) );
  XNOR2X1 U818 ( .A(n678), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n667), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n670), .B0(n672), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n671), .Y(n781) );
  XNOR2X1 U826 ( .A(n671), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule


module PE_0 ( rst_n, clk, inA, inB, inW, outC, outD );
  input [15:0] inA;
  input [39:0] inB;
  input [15:0] inW;
  output [39:0] outC;
  output [15:0] outD;
  input rst_n, clk;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N9, N8,
         N7, N6, N5, N4, N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23,
         N22, N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10,
         N1, n1;

  PE_0_DW_mult_tc_0 mult_971 ( .a(inA), .b(inW), .product({N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  PE_0_DW01_add_0 add_971 ( .A({n1, n1, n1, n1, n1, n1, n1, n1, n1, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), 
        .B(inB), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33}) );
  DFFRHQX1 outC_reg_39_ ( .D(N72), .CK(clk), .RN(rst_n), .Q(outC[39]) );
  DFFRHQX1 outC_reg_38_ ( .D(N71), .CK(clk), .RN(rst_n), .Q(outC[38]) );
  DFFRHQX1 outC_reg_37_ ( .D(N70), .CK(clk), .RN(rst_n), .Q(outC[37]) );
  DFFRHQX1 outC_reg_36_ ( .D(N69), .CK(clk), .RN(rst_n), .Q(outC[36]) );
  DFFRHQX1 outC_reg_35_ ( .D(N68), .CK(clk), .RN(rst_n), .Q(outC[35]) );
  DFFRHQX1 outC_reg_34_ ( .D(N67), .CK(clk), .RN(rst_n), .Q(outC[34]) );
  DFFRHQX1 outC_reg_33_ ( .D(N66), .CK(clk), .RN(rst_n), .Q(outC[33]) );
  DFFRHQX1 outC_reg_32_ ( .D(N65), .CK(clk), .RN(rst_n), .Q(outC[32]) );
  DFFRHQX1 outC_reg_31_ ( .D(N64), .CK(clk), .RN(rst_n), .Q(outC[31]) );
  DFFRHQX1 outC_reg_30_ ( .D(N63), .CK(clk), .RN(rst_n), .Q(outC[30]) );
  DFFRHQX1 outC_reg_29_ ( .D(N62), .CK(clk), .RN(rst_n), .Q(outC[29]) );
  DFFRHQX1 outC_reg_28_ ( .D(N61), .CK(clk), .RN(rst_n), .Q(outC[28]) );
  DFFRHQX1 outC_reg_27_ ( .D(N60), .CK(clk), .RN(rst_n), .Q(outC[27]) );
  DFFRHQX1 outC_reg_26_ ( .D(N59), .CK(clk), .RN(rst_n), .Q(outC[26]) );
  DFFRHQX1 outC_reg_25_ ( .D(N58), .CK(clk), .RN(rst_n), .Q(outC[25]) );
  DFFRHQX1 outC_reg_24_ ( .D(N57), .CK(clk), .RN(rst_n), .Q(outC[24]) );
  DFFRHQX1 outC_reg_23_ ( .D(N56), .CK(clk), .RN(rst_n), .Q(outC[23]) );
  DFFRHQX1 outC_reg_22_ ( .D(N55), .CK(clk), .RN(rst_n), .Q(outC[22]) );
  DFFRHQX1 outC_reg_21_ ( .D(N54), .CK(clk), .RN(rst_n), .Q(outC[21]) );
  DFFRHQX1 outC_reg_20_ ( .D(N53), .CK(clk), .RN(rst_n), .Q(outC[20]) );
  DFFRHQX1 outC_reg_19_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(outC[19]) );
  DFFRHQX1 outC_reg_18_ ( .D(N51), .CK(clk), .RN(rst_n), .Q(outC[18]) );
  DFFRHQX1 outC_reg_17_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(outC[17]) );
  DFFRHQX1 outC_reg_16_ ( .D(N49), .CK(clk), .RN(rst_n), .Q(outC[16]) );
  DFFRHQX1 outC_reg_15_ ( .D(N48), .CK(clk), .RN(rst_n), .Q(outC[15]) );
  DFFRHQX1 outC_reg_14_ ( .D(N47), .CK(clk), .RN(rst_n), .Q(outC[14]) );
  DFFRHQX1 outC_reg_13_ ( .D(N46), .CK(clk), .RN(rst_n), .Q(outC[13]) );
  DFFRHQX1 outC_reg_12_ ( .D(N45), .CK(clk), .RN(rst_n), .Q(outC[12]) );
  DFFRHQX1 outC_reg_11_ ( .D(N44), .CK(clk), .RN(rst_n), .Q(outC[11]) );
  DFFRHQX1 outC_reg_10_ ( .D(N43), .CK(clk), .RN(rst_n), .Q(outC[10]) );
  DFFRHQX1 outC_reg_9_ ( .D(N42), .CK(clk), .RN(rst_n), .Q(outC[9]) );
  DFFRHQX1 outC_reg_8_ ( .D(N41), .CK(clk), .RN(rst_n), .Q(outC[8]) );
  DFFRHQX1 outC_reg_7_ ( .D(N40), .CK(clk), .RN(rst_n), .Q(outC[7]) );
  DFFRHQX1 outC_reg_6_ ( .D(N39), .CK(clk), .RN(rst_n), .Q(outC[6]) );
  DFFRHQX1 outC_reg_5_ ( .D(N38), .CK(clk), .RN(rst_n), .Q(outC[5]) );
  DFFRHQX1 outC_reg_4_ ( .D(N37), .CK(clk), .RN(rst_n), .Q(outC[4]) );
  DFFRHQX1 outD_reg_14_ ( .D(inA[14]), .CK(clk), .RN(rst_n), .Q(outD[14]) );
  DFFRHQX1 outC_reg_3_ ( .D(N36), .CK(clk), .RN(rst_n), .Q(outC[3]) );
  DFFRHQX1 outC_reg_2_ ( .D(N35), .CK(clk), .RN(rst_n), .Q(outC[2]) );
  DFFRHQX1 outC_reg_1_ ( .D(N34), .CK(clk), .RN(rst_n), .Q(outC[1]) );
  DFFRHQX1 outC_reg_0_ ( .D(N33), .CK(clk), .RN(rst_n), .Q(outC[0]) );
  DFFRHQX1 outD_reg_15_ ( .D(inA[15]), .CK(clk), .RN(rst_n), .Q(outD[15]) );
  DFFRHQX1 outD_reg_12_ ( .D(inA[12]), .CK(clk), .RN(rst_n), .Q(outD[12]) );
  DFFRHQX1 outD_reg_10_ ( .D(inA[10]), .CK(clk), .RN(rst_n), .Q(outD[10]) );
  DFFRHQX1 outD_reg_8_ ( .D(inA[8]), .CK(clk), .RN(rst_n), .Q(outD[8]) );
  DFFRHQX1 outD_reg_13_ ( .D(inA[13]), .CK(clk), .RN(rst_n), .Q(outD[13]) );
  DFFRHQX1 outD_reg_11_ ( .D(inA[11]), .CK(clk), .RN(rst_n), .Q(outD[11]) );
  DFFRHQX1 outD_reg_6_ ( .D(inA[6]), .CK(clk), .RN(rst_n), .Q(outD[6]) );
  DFFRHQX1 outD_reg_4_ ( .D(inA[4]), .CK(clk), .RN(rst_n), .Q(outD[4]) );
  DFFRHQX1 outD_reg_2_ ( .D(inA[2]), .CK(clk), .RN(rst_n), .Q(outD[2]) );
  DFFRHQX1 outD_reg_9_ ( .D(inA[9]), .CK(clk), .RN(rst_n), .Q(outD[9]) );
  DFFRHQX1 outD_reg_7_ ( .D(inA[7]), .CK(clk), .RN(rst_n), .Q(outD[7]) );
  DFFRHQX1 outD_reg_5_ ( .D(inA[5]), .CK(clk), .RN(rst_n), .Q(outD[5]) );
  DFFRHQX1 outD_reg_0_ ( .D(inA[0]), .CK(clk), .RN(rst_n), .Q(outD[0]) );
  DFFRHQX1 outD_reg_3_ ( .D(inA[3]), .CK(clk), .RN(rst_n), .Q(outD[3]) );
  DFFRHQX1 outD_reg_1_ ( .D(inA[1]), .CK(clk), .RN(rst_n), .Q(outD[1]) );
  BUFX3 U3 ( .A(N32), .Y(n1) );
endmodule


module PE_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [39:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  XOR3X2 U1_39 ( .A(A[39]), .B(B[39]), .C(carry[39]), .Y(SUM[39]) );
  ADDFX2 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  ADDFX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  ADDFX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  ADDFX2 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFX2 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFX2 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFX2 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFX2 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  NOR2X1 U1 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  INVX1 U3 ( .A(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module PE_0_DW_mult_tc_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838;

  ADDFX2 U52 ( .A(n268), .B(n658), .CI(n52), .CO(n51), .S(product[30]) );
  ADDFX2 U53 ( .A(n83), .B(n82), .CI(n53), .CO(n52), .S(product[29]) );
  ADDFX2 U54 ( .A(n85), .B(n84), .CI(n54), .CO(n53), .S(product[28]) );
  ADDFX2 U55 ( .A(n90), .B(n86), .CI(n55), .CO(n54), .S(product[27]) );
  ADDFX2 U56 ( .A(n93), .B(n91), .CI(n56), .CO(n55), .S(product[26]) );
  ADDFX2 U57 ( .A(n94), .B(n98), .CI(n57), .CO(n56), .S(product[25]) );
  ADDFX2 U58 ( .A(n103), .B(n99), .CI(n58), .CO(n57), .S(product[24]) );
  ADDFX2 U59 ( .A(n104), .B(n110), .CI(n59), .CO(n58), .S(product[23]) );
  ADDFX2 U60 ( .A(n111), .B(n116), .CI(n60), .CO(n59), .S(product[22]) );
  ADDFX2 U61 ( .A(n117), .B(n124), .CI(n61), .CO(n60), .S(product[21]) );
  ADDFX2 U62 ( .A(n125), .B(n132), .CI(n62), .CO(n61), .S(product[20]) );
  ADDFX2 U63 ( .A(n142), .B(n133), .CI(n63), .CO(n62), .S(product[19]) );
  ADDFX2 U64 ( .A(n143), .B(n151), .CI(n64), .CO(n63), .S(product[18]) );
  ADDFX2 U65 ( .A(n152), .B(n162), .CI(n65), .CO(n64), .S(product[17]) );
  ADDFX2 U66 ( .A(n163), .B(n173), .CI(n66), .CO(n65), .S(product[16]) );
  ADDFX2 U67 ( .A(n174), .B(n184), .CI(n67), .CO(n66), .S(product[15]) );
  ADDFX2 U68 ( .A(n185), .B(n193), .CI(n68), .CO(n67), .S(product[14]) );
  ADDFX2 U69 ( .A(n194), .B(n203), .CI(n69), .CO(n68), .S(product[13]) );
  ADDFX2 U70 ( .A(n204), .B(n211), .CI(n70), .CO(n69), .S(product[12]) );
  ADDFX2 U71 ( .A(n212), .B(n219), .CI(n71), .CO(n70), .S(product[11]) );
  ADDFX2 U72 ( .A(n220), .B(n225), .CI(n72), .CO(n71), .S(product[10]) );
  ADDFX2 U73 ( .A(n226), .B(n232), .CI(n73), .CO(n72), .S(product[9]) );
  ADDFX2 U74 ( .A(n233), .B(n237), .CI(n74), .CO(n73), .S(product[8]) );
  ADDFX2 U75 ( .A(n238), .B(n242), .CI(n75), .CO(n74), .S(product[7]) );
  ADDFX2 U76 ( .A(n243), .B(n244), .CI(n76), .CO(n75), .S(product[6]) );
  ADDFX2 U77 ( .A(n245), .B(n248), .CI(n77), .CO(n76), .S(product[5]) );
  ADDFX2 U78 ( .A(n249), .B(n250), .CI(n78), .CO(n77), .S(product[4]) );
  ADDFX2 U79 ( .A(n251), .B(n266), .CI(n79), .CO(n78), .S(product[3]) );
  ADDFX2 U80 ( .A(n394), .B(n379), .CI(n80), .CO(n79), .S(product[2]) );
  ADDFX2 U83 ( .A(n269), .B(n657), .CI(n284), .CO(n83), .S(n84) );
  ADDFX2 U84 ( .A(n88), .B(n270), .CI(n89), .CO(n85), .S(n86) );
  CMPR42X1 U86 ( .A(n656), .B(n271), .C(n285), .D(n300), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U87 ( .A(n286), .B(n272), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U89 ( .A(n301), .B(n661), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFX2 U90 ( .A(n287), .B(n273), .CI(n315), .CO(n100), .S(n101) );
  CMPR42X1 U91 ( .A(n302), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFX2 U92 ( .A(n288), .B(n274), .CI(n108), .CO(n105), .S(n106) );
  CMPR42X1 U94 ( .A(n303), .B(n289), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U95 ( .A(n275), .B(n121), .C(n316), .D(n331), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U96 ( .A(n276), .B(n126), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U97 ( .A(n290), .B(n332), .C(n317), .D(n662), .ICI(n129), .S(n120), 
        .ICO(n118), .CO(n119) );
  CMPR42X1 U99 ( .A(n134), .B(n137), .C(n128), .D(n135), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U100 ( .A(n304), .B(n333), .C(n318), .D(n291), .ICI(n130), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFX2 U101 ( .A(n660), .B(n277), .CI(n348), .CO(n129), .S(n130) );
  CMPR42X1 U102 ( .A(n147), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U103 ( .A(n319), .B(n278), .C(n305), .D(n144), .ICI(n138), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFX2 U104 ( .A(n334), .B(n292), .CI(n140), .CO(n137), .S(n138) );
  CMPR42X1 U106 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U107 ( .A(n293), .B(n320), .C(n306), .D(n659), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U108 ( .A(n279), .B(n349), .C(n335), .D(n364), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U109 ( .A(n168), .B(n158), .C(n155), .D(n165), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U110 ( .A(n307), .B(n336), .C(n321), .D(n280), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U111 ( .A(n294), .B(n350), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CMPR42X1 U113 ( .A(n179), .B(n176), .C(n169), .D(n166), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U114 ( .A(n351), .B(n281), .C(n308), .D(n175), .ICI(n178), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U115 ( .A(n322), .B(n365), .C(n380), .D(n181), .ICI(n171), .S(n169), 
        .ICO(n167), .CO(n168) );
  CMPR42X1 U118 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U119 ( .A(n282), .B(n296), .C(n309), .D(n182), .ICI(n189), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U120 ( .A(n323), .B(n366), .C(n352), .D(n338), .ICI(n186), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U121 ( .A(n381), .B(n260), .CO(n181), .S(n182) );
  CMPR42X1 U122 ( .A(n353), .B(n191), .C(n196), .D(n188), .ICI(n192), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U123 ( .A(n367), .B(n324), .C(n339), .D(n200), .ICI(n198), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U124 ( .A(n283), .B(n382), .C(n297), .D(n310), .ICI(n195), .S(n191), 
        .ICO(n189), .CO(n190) );
  CMPR42X1 U125 ( .A(n205), .B(n208), .C(n206), .D(n197), .ICI(n202), .S(n194), 
        .ICO(n192), .CO(n193) );
  CMPR42X1 U126 ( .A(n354), .B(n311), .C(n340), .D(n201), .ICI(n199), .S(n197), 
        .ICO(n195), .CO(n196) );
  ADDFX2 U127 ( .A(n368), .B(n325), .CI(n298), .CO(n198), .S(n199) );
  ADDHXL U128 ( .A(n383), .B(n261), .CO(n200), .S(n201) );
  CMPR42X1 U129 ( .A(n341), .B(n213), .C(n214), .D(n207), .ICI(n210), .S(n204), 
        .ICO(n202), .CO(n203) );
  CMPR42X1 U130 ( .A(n369), .B(n326), .C(n355), .D(n216), .ICI(n209), .S(n207), 
        .ICO(n205), .CO(n206) );
  ADDFX2 U131 ( .A(n384), .B(n299), .CI(n312), .CO(n208), .S(n209) );
  CMPR42X1 U132 ( .A(n327), .B(n217), .C(n218), .D(n222), .ICI(n215), .S(n212), 
        .ICO(n210), .CO(n211) );
  CMPR42X1 U133 ( .A(n342), .B(n370), .C(n356), .D(n313), .ICI(n221), .S(n215), 
        .ICO(n213), .CO(n214) );
  CMPR42X1 U135 ( .A(n371), .B(n357), .C(n227), .D(n224), .ICI(n223), .S(n220), 
        .ICO(n218), .CO(n219) );
  CMPR42X1 U136 ( .A(n314), .B(n386), .C(n328), .D(n343), .ICI(n229), .S(n223), 
        .ICO(n221), .CO(n222) );
  CMPR42X1 U137 ( .A(n372), .B(n230), .C(n234), .D(n231), .ICI(n228), .S(n226), 
        .ICO(n224), .CO(n225) );
  ADDFX2 U138 ( .A(n329), .B(n344), .CI(n358), .CO(n227), .S(n228) );
  CMPR42X1 U140 ( .A(n373), .B(n359), .C(n239), .D(n236), .ICI(n235), .S(n233), 
        .ICO(n231), .CO(n232) );
  ADDFX2 U141 ( .A(n388), .B(n330), .CI(n345), .CO(n234), .S(n235) );
  CMPR42X1 U142 ( .A(n374), .B(n346), .C(n360), .D(n240), .ICI(n241), .S(n238), 
        .ICO(n236), .CO(n237) );
  CMPR42X1 U144 ( .A(n347), .B(n390), .C(n361), .D(n375), .ICI(n246), .S(n243), 
        .ICO(n241), .CO(n242) );
  ADDFX2 U145 ( .A(n362), .B(n376), .CI(n247), .CO(n244), .S(n245) );
  ADDHXL U146 ( .A(n391), .B(n265), .CO(n246), .S(n247) );
  ADDFX2 U147 ( .A(n392), .B(n363), .CI(n377), .CO(n248), .S(n249) );
  CMPR22X1 U486 ( .A(n267), .B(n395), .CO(n80), .S(product[1]) );
  CMPR22X1 U487 ( .A(n387), .B(n263), .CO(n229), .S(n230) );
  CMPR22X1 U488 ( .A(n385), .B(n262), .CO(n216), .S(n217) );
  CMPR22X1 U489 ( .A(n393), .B(n378), .CO(n250), .S(n251) );
  CMPR22X1 U490 ( .A(n389), .B(n264), .CO(n239), .S(n240) );
  INVX1 U491 ( .A(n160), .Y(n659) );
  INVX1 U492 ( .A(n121), .Y(n662) );
  INVX1 U493 ( .A(n96), .Y(n656) );
  INVX1 U494 ( .A(n82), .Y(n658) );
  CLKINVX3 U495 ( .A(n709), .Y(n685) );
  CLKINVX3 U496 ( .A(n649), .Y(n683) );
  INVX1 U497 ( .A(n648), .Y(n686) );
  CLKINVX3 U498 ( .A(n651), .Y(n677) );
  CLKINVX3 U499 ( .A(n650), .Y(n680) );
  CLKINVX3 U500 ( .A(n652), .Y(n674) );
  CLKINVX3 U501 ( .A(n647), .Y(n663) );
  CLKINVX3 U502 ( .A(n653), .Y(n671) );
  CLKINVX3 U503 ( .A(n654), .Y(n668) );
  INVX1 U504 ( .A(n710), .Y(n684) );
  INVX1 U505 ( .A(n712), .Y(n682) );
  INVX1 U506 ( .A(n655), .Y(n665) );
  INVX1 U507 ( .A(n728), .Y(n681) );
  INVX1 U508 ( .A(n730), .Y(n679) );
  INVX1 U509 ( .A(n140), .Y(n660) );
  INVX1 U510 ( .A(n746), .Y(n678) );
  INVX1 U511 ( .A(n764), .Y(n675) );
  INVX1 U512 ( .A(n766), .Y(n673) );
  INVX1 U513 ( .A(n748), .Y(n676) );
  INVX1 U514 ( .A(n108), .Y(n661) );
  INVX1 U515 ( .A(n782), .Y(n672) );
  INVX1 U516 ( .A(n784), .Y(n670) );
  INVX1 U517 ( .A(n798), .Y(n669) );
  INVX1 U518 ( .A(n800), .Y(n667) );
  INVX1 U519 ( .A(n88), .Y(n657) );
  INVX1 U520 ( .A(n814), .Y(n666) );
  INVX1 U521 ( .A(n816), .Y(n664) );
  XOR2X2 U522 ( .A(a[4]), .B(n683), .Y(n728) );
  XOR2X2 U523 ( .A(a[2]), .B(n686), .Y(n710) );
  BUFX3 U524 ( .A(a[3]), .Y(n649) );
  BUFX3 U525 ( .A(a[1]), .Y(n648) );
  XOR2X2 U526 ( .A(a[6]), .B(n680), .Y(n746) );
  XOR2X2 U527 ( .A(a[8]), .B(n677), .Y(n764) );
  CLKINVX3 U528 ( .A(a[0]), .Y(n687) );
  BUFX3 U529 ( .A(a[7]), .Y(n651) );
  BUFX3 U530 ( .A(a[5]), .Y(n650) );
  BUFX3 U531 ( .A(a[9]), .Y(n652) );
  BUFX3 U532 ( .A(b[0]), .Y(n647) );
  XOR2X2 U533 ( .A(a[10]), .B(n674), .Y(n782) );
  XOR2X2 U534 ( .A(a[12]), .B(n671), .Y(n798) );
  BUFX3 U535 ( .A(a[11]), .Y(n653) );
  BUFX3 U536 ( .A(a[13]), .Y(n654) );
  XOR2X2 U537 ( .A(a[14]), .B(n668), .Y(n814) );
  BUFX3 U538 ( .A(a[15]), .Y(n655) );
  NAND2X4 U539 ( .A(n814), .B(n830), .Y(n816) );
  NAND2X4 U540 ( .A(n746), .B(n833), .Y(n748) );
  NAND2X4 U541 ( .A(n798), .B(n834), .Y(n800) );
  NAND2X4 U542 ( .A(n710), .B(n835), .Y(n712) );
  NAND2X4 U543 ( .A(n728), .B(n836), .Y(n730) );
  NAND2X4 U544 ( .A(n782), .B(n837), .Y(n784) );
  NAND2X4 U545 ( .A(n764), .B(n838), .Y(n766) );
  INVX1 U546 ( .A(n51), .Y(product[31]) );
  NOR2X1 U547 ( .A(n687), .B(n663), .Y(product[0]) );
  AOI22X1 U548 ( .A0(n688), .A1(n670), .B0(n672), .B1(n689), .Y(n96) );
  AOI22X1 U549 ( .A0(n690), .A1(n667), .B0(n669), .B1(n691), .Y(n88) );
  AOI22X1 U550 ( .A0(n692), .A1(n664), .B0(n666), .B1(n693), .Y(n82) );
  OAI22X1 U551 ( .A0(n647), .A1(n685), .B0(n694), .B1(n687), .Y(n395) );
  OAI22X1 U552 ( .A0(n694), .A1(n685), .B0(n695), .B1(n687), .Y(n394) );
  XNOR2X1 U553 ( .A(b[1]), .B(n648), .Y(n694) );
  OAI22X1 U554 ( .A0(n695), .A1(n685), .B0(n696), .B1(n687), .Y(n393) );
  XNOR2X1 U555 ( .A(b[2]), .B(n648), .Y(n695) );
  OAI22X1 U556 ( .A0(n696), .A1(n685), .B0(n697), .B1(n687), .Y(n392) );
  XNOR2X1 U557 ( .A(b[3]), .B(n648), .Y(n696) );
  OAI22X1 U558 ( .A0(n697), .A1(n685), .B0(n698), .B1(n687), .Y(n391) );
  XNOR2X1 U559 ( .A(b[4]), .B(n648), .Y(n697) );
  OAI22X1 U560 ( .A0(n698), .A1(n685), .B0(n699), .B1(n687), .Y(n390) );
  XNOR2X1 U561 ( .A(b[5]), .B(n648), .Y(n698) );
  OAI22X1 U562 ( .A0(n699), .A1(n685), .B0(n700), .B1(n687), .Y(n389) );
  XNOR2X1 U563 ( .A(b[6]), .B(n648), .Y(n699) );
  OAI22X1 U564 ( .A0(n700), .A1(n685), .B0(n701), .B1(n687), .Y(n388) );
  XNOR2X1 U565 ( .A(b[7]), .B(n648), .Y(n700) );
  OAI22X1 U566 ( .A0(n701), .A1(n685), .B0(n702), .B1(n687), .Y(n387) );
  XNOR2X1 U567 ( .A(b[8]), .B(n648), .Y(n701) );
  OAI22X1 U568 ( .A0(n702), .A1(n685), .B0(n703), .B1(n687), .Y(n386) );
  XNOR2X1 U569 ( .A(b[9]), .B(n648), .Y(n702) );
  OAI22X1 U570 ( .A0(n703), .A1(n685), .B0(n704), .B1(n687), .Y(n385) );
  XNOR2X1 U571 ( .A(b[10]), .B(n648), .Y(n703) );
  OAI22X1 U572 ( .A0(n704), .A1(n685), .B0(n705), .B1(n687), .Y(n384) );
  XNOR2X1 U573 ( .A(b[11]), .B(n648), .Y(n704) );
  OAI22X1 U574 ( .A0(n705), .A1(n685), .B0(n706), .B1(n687), .Y(n383) );
  XNOR2X1 U575 ( .A(b[12]), .B(n648), .Y(n705) );
  OAI22X1 U576 ( .A0(n706), .A1(n685), .B0(n707), .B1(n687), .Y(n382) );
  XNOR2X1 U577 ( .A(b[13]), .B(n648), .Y(n706) );
  OAI2BB2X1 U578 ( .B0(n707), .B1(n685), .A0N(n708), .A1N(a[0]), .Y(n381) );
  XNOR2X1 U579 ( .A(b[14]), .B(n648), .Y(n707) );
  AOI22X1 U580 ( .A0(a[0]), .A1(n708), .B0(n709), .B1(n708), .Y(n380) );
  XNOR2X1 U581 ( .A(b[15]), .B(n686), .Y(n708) );
  NOR2X1 U582 ( .A(n710), .B(n663), .Y(n379) );
  OAI22X1 U583 ( .A0(n711), .A1(n712), .B0(n710), .B1(n713), .Y(n378) );
  XNOR2X1 U584 ( .A(n649), .B(n647), .Y(n711) );
  OAI22X1 U585 ( .A0(n713), .A1(n712), .B0(n710), .B1(n714), .Y(n377) );
  XNOR2X1 U586 ( .A(b[1]), .B(n649), .Y(n713) );
  OAI22X1 U587 ( .A0(n714), .A1(n712), .B0(n710), .B1(n715), .Y(n376) );
  XNOR2X1 U588 ( .A(b[2]), .B(n649), .Y(n714) );
  OAI22X1 U589 ( .A0(n715), .A1(n712), .B0(n710), .B1(n716), .Y(n375) );
  XNOR2X1 U590 ( .A(b[3]), .B(n649), .Y(n715) );
  OAI22X1 U591 ( .A0(n716), .A1(n712), .B0(n710), .B1(n717), .Y(n374) );
  XNOR2X1 U592 ( .A(b[4]), .B(n649), .Y(n716) );
  OAI22X1 U593 ( .A0(n717), .A1(n712), .B0(n710), .B1(n718), .Y(n373) );
  XNOR2X1 U594 ( .A(b[5]), .B(n649), .Y(n717) );
  OAI22X1 U595 ( .A0(n718), .A1(n712), .B0(n710), .B1(n719), .Y(n372) );
  XNOR2X1 U596 ( .A(b[6]), .B(n649), .Y(n718) );
  OAI22X1 U597 ( .A0(n719), .A1(n712), .B0(n710), .B1(n720), .Y(n371) );
  XNOR2X1 U598 ( .A(b[7]), .B(n649), .Y(n719) );
  OAI22X1 U599 ( .A0(n720), .A1(n712), .B0(n710), .B1(n721), .Y(n370) );
  XNOR2X1 U600 ( .A(b[8]), .B(n649), .Y(n720) );
  OAI22X1 U601 ( .A0(n721), .A1(n712), .B0(n710), .B1(n722), .Y(n369) );
  XNOR2X1 U602 ( .A(b[9]), .B(n649), .Y(n721) );
  OAI22X1 U603 ( .A0(n722), .A1(n712), .B0(n710), .B1(n723), .Y(n368) );
  XNOR2X1 U604 ( .A(b[10]), .B(n649), .Y(n722) );
  OAI22X1 U605 ( .A0(n723), .A1(n712), .B0(n710), .B1(n724), .Y(n367) );
  XNOR2X1 U606 ( .A(b[11]), .B(n649), .Y(n723) );
  OAI22X1 U607 ( .A0(n724), .A1(n712), .B0(n710), .B1(n725), .Y(n366) );
  XNOR2X1 U608 ( .A(b[12]), .B(n649), .Y(n724) );
  OAI2BB2X1 U609 ( .B0(n725), .B1(n712), .A0N(n684), .A1N(n726), .Y(n365) );
  XNOR2X1 U610 ( .A(b[13]), .B(n649), .Y(n725) );
  AOI22X1 U611 ( .A0(n727), .A1(n684), .B0(n682), .B1(n727), .Y(n364) );
  NOR2X1 U612 ( .A(n728), .B(n663), .Y(n363) );
  OAI22X1 U613 ( .A0(n729), .A1(n730), .B0(n728), .B1(n731), .Y(n362) );
  XNOR2X1 U614 ( .A(n650), .B(n647), .Y(n729) );
  OAI22X1 U615 ( .A0(n731), .A1(n730), .B0(n728), .B1(n732), .Y(n361) );
  XNOR2X1 U616 ( .A(b[1]), .B(n650), .Y(n731) );
  OAI22X1 U617 ( .A0(n732), .A1(n730), .B0(n728), .B1(n733), .Y(n360) );
  XNOR2X1 U618 ( .A(b[2]), .B(n650), .Y(n732) );
  OAI22X1 U619 ( .A0(n733), .A1(n730), .B0(n728), .B1(n734), .Y(n359) );
  XNOR2X1 U620 ( .A(b[3]), .B(n650), .Y(n733) );
  OAI22X1 U621 ( .A0(n734), .A1(n730), .B0(n728), .B1(n735), .Y(n358) );
  XNOR2X1 U622 ( .A(b[4]), .B(n650), .Y(n734) );
  OAI22X1 U623 ( .A0(n735), .A1(n730), .B0(n728), .B1(n736), .Y(n357) );
  XNOR2X1 U624 ( .A(b[5]), .B(n650), .Y(n735) );
  OAI22X1 U625 ( .A0(n736), .A1(n730), .B0(n728), .B1(n737), .Y(n356) );
  XNOR2X1 U626 ( .A(b[6]), .B(n650), .Y(n736) );
  OAI22X1 U627 ( .A0(n737), .A1(n730), .B0(n728), .B1(n738), .Y(n355) );
  XNOR2X1 U628 ( .A(b[7]), .B(n650), .Y(n737) );
  OAI22X1 U629 ( .A0(n738), .A1(n730), .B0(n728), .B1(n739), .Y(n354) );
  XNOR2X1 U630 ( .A(b[8]), .B(n650), .Y(n738) );
  OAI22X1 U631 ( .A0(n739), .A1(n730), .B0(n728), .B1(n740), .Y(n353) );
  XNOR2X1 U632 ( .A(b[9]), .B(n650), .Y(n739) );
  OAI22X1 U633 ( .A0(n740), .A1(n730), .B0(n728), .B1(n741), .Y(n352) );
  XNOR2X1 U634 ( .A(b[10]), .B(n650), .Y(n740) );
  OAI22X1 U635 ( .A0(n741), .A1(n730), .B0(n728), .B1(n742), .Y(n351) );
  XNOR2X1 U636 ( .A(b[11]), .B(n650), .Y(n741) );
  OAI22X1 U637 ( .A0(n742), .A1(n730), .B0(n728), .B1(n743), .Y(n350) );
  XNOR2X1 U638 ( .A(b[12]), .B(n650), .Y(n742) );
  OAI2BB2X1 U639 ( .B0(n743), .B1(n730), .A0N(n681), .A1N(n744), .Y(n349) );
  XNOR2X1 U640 ( .A(b[13]), .B(n650), .Y(n743) );
  AOI22X1 U641 ( .A0(n745), .A1(n681), .B0(n679), .B1(n745), .Y(n348) );
  NOR2X1 U642 ( .A(n746), .B(n663), .Y(n347) );
  OAI22X1 U643 ( .A0(n747), .A1(n748), .B0(n746), .B1(n749), .Y(n346) );
  XNOR2X1 U644 ( .A(n651), .B(n647), .Y(n747) );
  OAI22X1 U645 ( .A0(n749), .A1(n748), .B0(n746), .B1(n750), .Y(n345) );
  XNOR2X1 U646 ( .A(b[1]), .B(n651), .Y(n749) );
  OAI22X1 U647 ( .A0(n750), .A1(n748), .B0(n746), .B1(n751), .Y(n344) );
  XNOR2X1 U648 ( .A(b[2]), .B(n651), .Y(n750) );
  OAI22X1 U649 ( .A0(n751), .A1(n748), .B0(n746), .B1(n752), .Y(n343) );
  XNOR2X1 U650 ( .A(b[3]), .B(n651), .Y(n751) );
  OAI22X1 U651 ( .A0(n752), .A1(n748), .B0(n746), .B1(n753), .Y(n342) );
  XNOR2X1 U652 ( .A(b[4]), .B(n651), .Y(n752) );
  OAI22X1 U653 ( .A0(n753), .A1(n748), .B0(n746), .B1(n754), .Y(n341) );
  XNOR2X1 U654 ( .A(b[5]), .B(n651), .Y(n753) );
  OAI22X1 U655 ( .A0(n754), .A1(n748), .B0(n746), .B1(n755), .Y(n340) );
  XNOR2X1 U656 ( .A(b[6]), .B(n651), .Y(n754) );
  OAI22X1 U657 ( .A0(n755), .A1(n748), .B0(n746), .B1(n756), .Y(n339) );
  XNOR2X1 U658 ( .A(b[7]), .B(n651), .Y(n755) );
  OAI22X1 U659 ( .A0(n756), .A1(n748), .B0(n746), .B1(n757), .Y(n338) );
  XNOR2X1 U660 ( .A(b[8]), .B(n651), .Y(n756) );
  OAI22X1 U661 ( .A0(n758), .A1(n748), .B0(n746), .B1(n759), .Y(n336) );
  OAI22X1 U662 ( .A0(n759), .A1(n748), .B0(n746), .B1(n760), .Y(n335) );
  XNOR2X1 U663 ( .A(b[11]), .B(n651), .Y(n759) );
  OAI22X1 U664 ( .A0(n760), .A1(n748), .B0(n746), .B1(n761), .Y(n334) );
  XNOR2X1 U665 ( .A(b[12]), .B(n651), .Y(n760) );
  OAI22X1 U666 ( .A0(n761), .A1(n748), .B0(n746), .B1(n762), .Y(n333) );
  XNOR2X1 U667 ( .A(b[13]), .B(n651), .Y(n761) );
  OAI2BB2X1 U668 ( .B0(n762), .B1(n748), .A0N(n678), .A1N(n763), .Y(n332) );
  XNOR2X1 U669 ( .A(b[14]), .B(n651), .Y(n762) );
  AOI22X1 U670 ( .A0(n763), .A1(n678), .B0(n676), .B1(n763), .Y(n331) );
  XNOR2X1 U671 ( .A(b[15]), .B(n677), .Y(n763) );
  NOR2X1 U672 ( .A(n764), .B(n663), .Y(n330) );
  OAI22X1 U673 ( .A0(n765), .A1(n766), .B0(n764), .B1(n767), .Y(n329) );
  XNOR2X1 U674 ( .A(n652), .B(n647), .Y(n765) );
  OAI22X1 U675 ( .A0(n767), .A1(n766), .B0(n764), .B1(n768), .Y(n328) );
  XNOR2X1 U676 ( .A(b[1]), .B(n652), .Y(n767) );
  OAI22X1 U677 ( .A0(n768), .A1(n766), .B0(n764), .B1(n769), .Y(n327) );
  XNOR2X1 U678 ( .A(b[2]), .B(n652), .Y(n768) );
  OAI22X1 U679 ( .A0(n769), .A1(n766), .B0(n764), .B1(n770), .Y(n326) );
  XNOR2X1 U680 ( .A(b[3]), .B(n652), .Y(n769) );
  OAI22X1 U681 ( .A0(n770), .A1(n766), .B0(n764), .B1(n771), .Y(n325) );
  XNOR2X1 U682 ( .A(b[4]), .B(n652), .Y(n770) );
  OAI22X1 U683 ( .A0(n771), .A1(n766), .B0(n764), .B1(n772), .Y(n324) );
  XNOR2X1 U684 ( .A(b[5]), .B(n652), .Y(n771) );
  OAI22X1 U685 ( .A0(n772), .A1(n766), .B0(n764), .B1(n773), .Y(n323) );
  XNOR2X1 U686 ( .A(b[6]), .B(n652), .Y(n772) );
  OAI22X1 U687 ( .A0(n773), .A1(n766), .B0(n764), .B1(n774), .Y(n322) );
  XNOR2X1 U688 ( .A(b[7]), .B(n652), .Y(n773) );
  OAI22X1 U689 ( .A0(n774), .A1(n766), .B0(n764), .B1(n775), .Y(n321) );
  XNOR2X1 U690 ( .A(b[8]), .B(n652), .Y(n774) );
  OAI22X1 U691 ( .A0(n775), .A1(n766), .B0(n764), .B1(n776), .Y(n320) );
  XNOR2X1 U692 ( .A(b[9]), .B(n652), .Y(n775) );
  OAI22X1 U693 ( .A0(n776), .A1(n766), .B0(n764), .B1(n777), .Y(n319) );
  XNOR2X1 U694 ( .A(b[10]), .B(n652), .Y(n776) );
  OAI22X1 U695 ( .A0(n777), .A1(n766), .B0(n764), .B1(n778), .Y(n318) );
  XNOR2X1 U696 ( .A(b[11]), .B(n652), .Y(n777) );
  OAI22X1 U697 ( .A0(n778), .A1(n766), .B0(n764), .B1(n779), .Y(n317) );
  XNOR2X1 U698 ( .A(b[12]), .B(n652), .Y(n778) );
  OAI2BB2X1 U699 ( .B0(n779), .B1(n766), .A0N(n675), .A1N(n780), .Y(n316) );
  XNOR2X1 U700 ( .A(b[13]), .B(n652), .Y(n779) );
  AOI22X1 U701 ( .A0(n781), .A1(n675), .B0(n673), .B1(n781), .Y(n315) );
  NOR2X1 U702 ( .A(n782), .B(n663), .Y(n314) );
  OAI22X1 U703 ( .A0(n783), .A1(n784), .B0(n782), .B1(n785), .Y(n313) );
  XNOR2X1 U704 ( .A(n653), .B(n647), .Y(n783) );
  OAI22X1 U705 ( .A0(n785), .A1(n784), .B0(n782), .B1(n786), .Y(n312) );
  XNOR2X1 U706 ( .A(b[1]), .B(n653), .Y(n785) );
  OAI22X1 U707 ( .A0(n786), .A1(n784), .B0(n782), .B1(n787), .Y(n311) );
  XNOR2X1 U708 ( .A(b[2]), .B(n653), .Y(n786) );
  OAI22X1 U709 ( .A0(n787), .A1(n784), .B0(n782), .B1(n788), .Y(n310) );
  XNOR2X1 U710 ( .A(b[3]), .B(n653), .Y(n787) );
  OAI22X1 U711 ( .A0(n788), .A1(n784), .B0(n782), .B1(n789), .Y(n309) );
  XNOR2X1 U712 ( .A(b[4]), .B(n653), .Y(n788) );
  OAI22X1 U713 ( .A0(n789), .A1(n784), .B0(n782), .B1(n790), .Y(n308) );
  XNOR2X1 U714 ( .A(b[5]), .B(n653), .Y(n789) );
  OAI22X1 U715 ( .A0(n790), .A1(n784), .B0(n782), .B1(n791), .Y(n307) );
  XNOR2X1 U716 ( .A(b[6]), .B(n653), .Y(n790) );
  OAI22X1 U717 ( .A0(n791), .A1(n784), .B0(n782), .B1(n792), .Y(n306) );
  XNOR2X1 U718 ( .A(b[7]), .B(n653), .Y(n791) );
  OAI22X1 U719 ( .A0(n792), .A1(n784), .B0(n782), .B1(n793), .Y(n305) );
  XNOR2X1 U720 ( .A(b[8]), .B(n653), .Y(n792) );
  OAI22X1 U721 ( .A0(n793), .A1(n784), .B0(n782), .B1(n794), .Y(n304) );
  XNOR2X1 U722 ( .A(b[9]), .B(n653), .Y(n793) );
  OAI22X1 U723 ( .A0(n795), .A1(n784), .B0(n782), .B1(n796), .Y(n303) );
  OAI22X1 U724 ( .A0(n796), .A1(n784), .B0(n782), .B1(n797), .Y(n302) );
  XNOR2X1 U725 ( .A(b[12]), .B(n653), .Y(n796) );
  OAI2BB2X1 U726 ( .B0(n797), .B1(n784), .A0N(n672), .A1N(n688), .Y(n301) );
  XOR2X1 U727 ( .A(b[14]), .B(n653), .Y(n688) );
  XNOR2X1 U728 ( .A(b[13]), .B(n653), .Y(n797) );
  AOI22X1 U729 ( .A0(n689), .A1(n672), .B0(n670), .B1(n689), .Y(n300) );
  XNOR2X1 U730 ( .A(b[15]), .B(n671), .Y(n689) );
  NOR2X1 U731 ( .A(n798), .B(n663), .Y(n299) );
  OAI22X1 U732 ( .A0(n799), .A1(n800), .B0(n798), .B1(n801), .Y(n298) );
  XNOR2X1 U733 ( .A(n654), .B(n647), .Y(n799) );
  OAI22X1 U734 ( .A0(n801), .A1(n800), .B0(n798), .B1(n802), .Y(n297) );
  XNOR2X1 U735 ( .A(b[1]), .B(n654), .Y(n801) );
  OAI22X1 U736 ( .A0(n802), .A1(n800), .B0(n798), .B1(n803), .Y(n296) );
  XNOR2X1 U737 ( .A(b[2]), .B(n654), .Y(n802) );
  OAI22X1 U738 ( .A0(n804), .A1(n800), .B0(n798), .B1(n805), .Y(n294) );
  OAI22X1 U739 ( .A0(n805), .A1(n800), .B0(n798), .B1(n806), .Y(n293) );
  XNOR2X1 U740 ( .A(b[5]), .B(n654), .Y(n805) );
  OAI22X1 U741 ( .A0(n806), .A1(n800), .B0(n798), .B1(n807), .Y(n292) );
  XNOR2X1 U742 ( .A(b[6]), .B(n654), .Y(n806) );
  OAI22X1 U743 ( .A0(n807), .A1(n800), .B0(n798), .B1(n808), .Y(n291) );
  XNOR2X1 U744 ( .A(b[7]), .B(n654), .Y(n807) );
  OAI22X1 U745 ( .A0(n808), .A1(n800), .B0(n798), .B1(n809), .Y(n290) );
  XNOR2X1 U746 ( .A(b[8]), .B(n654), .Y(n808) );
  OAI22X1 U747 ( .A0(n809), .A1(n800), .B0(n798), .B1(n810), .Y(n289) );
  XNOR2X1 U748 ( .A(b[9]), .B(n654), .Y(n809) );
  OAI22X1 U749 ( .A0(n810), .A1(n800), .B0(n798), .B1(n811), .Y(n288) );
  XNOR2X1 U750 ( .A(b[10]), .B(n654), .Y(n810) );
  OAI22X1 U751 ( .A0(n811), .A1(n800), .B0(n798), .B1(n812), .Y(n287) );
  XNOR2X1 U752 ( .A(b[11]), .B(n654), .Y(n811) );
  OAI22X1 U753 ( .A0(n812), .A1(n800), .B0(n798), .B1(n813), .Y(n286) );
  XNOR2X1 U754 ( .A(b[12]), .B(n654), .Y(n812) );
  OAI2BB2X1 U755 ( .B0(n813), .B1(n800), .A0N(n669), .A1N(n690), .Y(n285) );
  XOR2X1 U756 ( .A(b[14]), .B(n654), .Y(n690) );
  XNOR2X1 U757 ( .A(b[13]), .B(n654), .Y(n813) );
  AOI22X1 U758 ( .A0(n691), .A1(n669), .B0(n667), .B1(n691), .Y(n284) );
  XNOR2X1 U759 ( .A(b[15]), .B(n668), .Y(n691) );
  NOR2X1 U760 ( .A(n814), .B(n663), .Y(n283) );
  OAI22X1 U761 ( .A0(n815), .A1(n816), .B0(n814), .B1(n817), .Y(n282) );
  XNOR2X1 U762 ( .A(n655), .B(n647), .Y(n815) );
  OAI22X1 U763 ( .A0(n817), .A1(n816), .B0(n814), .B1(n818), .Y(n281) );
  XNOR2X1 U764 ( .A(b[1]), .B(n655), .Y(n817) );
  OAI22X1 U765 ( .A0(n818), .A1(n816), .B0(n814), .B1(n819), .Y(n280) );
  XNOR2X1 U766 ( .A(b[2]), .B(n655), .Y(n818) );
  OAI22X1 U767 ( .A0(n819), .A1(n816), .B0(n814), .B1(n820), .Y(n279) );
  XNOR2X1 U768 ( .A(b[3]), .B(n655), .Y(n819) );
  OAI22X1 U769 ( .A0(n820), .A1(n816), .B0(n814), .B1(n821), .Y(n278) );
  XNOR2X1 U770 ( .A(b[4]), .B(n655), .Y(n820) );
  OAI22X1 U771 ( .A0(n821), .A1(n816), .B0(n814), .B1(n822), .Y(n277) );
  XNOR2X1 U772 ( .A(b[5]), .B(n655), .Y(n821) );
  OAI22X1 U773 ( .A0(n822), .A1(n816), .B0(n814), .B1(n823), .Y(n276) );
  XNOR2X1 U774 ( .A(b[6]), .B(n655), .Y(n822) );
  OAI22X1 U775 ( .A0(n823), .A1(n816), .B0(n814), .B1(n824), .Y(n275) );
  XNOR2X1 U776 ( .A(b[7]), .B(n655), .Y(n823) );
  OAI22X1 U777 ( .A0(n824), .A1(n816), .B0(n814), .B1(n825), .Y(n274) );
  XNOR2X1 U778 ( .A(b[8]), .B(n655), .Y(n824) );
  OAI22X1 U779 ( .A0(n825), .A1(n816), .B0(n814), .B1(n826), .Y(n273) );
  XNOR2X1 U780 ( .A(b[9]), .B(n655), .Y(n825) );
  OAI22X1 U781 ( .A0(n826), .A1(n816), .B0(n814), .B1(n827), .Y(n272) );
  XNOR2X1 U782 ( .A(b[10]), .B(n655), .Y(n826) );
  OAI22X1 U783 ( .A0(n827), .A1(n816), .B0(n814), .B1(n828), .Y(n271) );
  XNOR2X1 U784 ( .A(b[11]), .B(n655), .Y(n827) );
  OAI22X1 U785 ( .A0(n828), .A1(n816), .B0(n814), .B1(n829), .Y(n270) );
  XNOR2X1 U786 ( .A(b[12]), .B(n655), .Y(n828) );
  OAI2BB2X1 U787 ( .B0(n829), .B1(n816), .A0N(n666), .A1N(n692), .Y(n269) );
  XOR2X1 U788 ( .A(b[14]), .B(n655), .Y(n692) );
  XNOR2X1 U789 ( .A(b[13]), .B(n655), .Y(n829) );
  AOI22X1 U790 ( .A0(n693), .A1(n666), .B0(n664), .B1(n693), .Y(n268) );
  XNOR2X1 U791 ( .A(b[15]), .B(n665), .Y(n693) );
  OAI21XL U792 ( .A0(n647), .A1(n686), .B0(n685), .Y(n267) );
  NOR2X1 U793 ( .A(n686), .B(a[0]), .Y(n709) );
  OAI32X1 U794 ( .A0(n683), .A1(n647), .A2(n710), .B0(n683), .B1(n712), .Y(
        n266) );
  OAI32X1 U795 ( .A0(n680), .A1(n647), .A2(n728), .B0(n680), .B1(n730), .Y(
        n265) );
  OAI32X1 U796 ( .A0(n677), .A1(n647), .A2(n746), .B0(n677), .B1(n748), .Y(
        n264) );
  OAI32X1 U797 ( .A0(n674), .A1(n647), .A2(n764), .B0(n674), .B1(n766), .Y(
        n263) );
  OAI32X1 U798 ( .A0(n671), .A1(n647), .A2(n782), .B0(n671), .B1(n784), .Y(
        n262) );
  OAI32X1 U799 ( .A0(n668), .A1(n647), .A2(n798), .B0(n668), .B1(n800), .Y(
        n261) );
  OAI32X1 U800 ( .A0(n665), .A1(n647), .A2(n814), .B0(n665), .B1(n816), .Y(
        n260) );
  XNOR2X1 U801 ( .A(n665), .B(a[14]), .Y(n830) );
  XNOR2X1 U802 ( .A(n831), .B(n832), .Y(n171) );
  OR2X1 U803 ( .A(n831), .B(n832), .Y(n170) );
  OAI22X1 U804 ( .A0(n757), .A1(n748), .B0(n746), .B1(n758), .Y(n832) );
  XNOR2X1 U805 ( .A(b[10]), .B(n651), .Y(n758) );
  XNOR2X1 U806 ( .A(n677), .B(a[6]), .Y(n833) );
  XNOR2X1 U807 ( .A(b[9]), .B(n651), .Y(n757) );
  OAI22X1 U808 ( .A0(n803), .A1(n800), .B0(n798), .B1(n804), .Y(n831) );
  XNOR2X1 U809 ( .A(b[4]), .B(n654), .Y(n804) );
  XNOR2X1 U810 ( .A(n668), .B(a[12]), .Y(n834) );
  XNOR2X1 U811 ( .A(b[3]), .B(n654), .Y(n803) );
  AOI22X1 U812 ( .A0(n726), .A1(n682), .B0(n684), .B1(n727), .Y(n160) );
  XNOR2X1 U813 ( .A(b[15]), .B(n683), .Y(n727) );
  XNOR2X1 U814 ( .A(n683), .B(a[2]), .Y(n835) );
  XOR2X1 U815 ( .A(b[14]), .B(n649), .Y(n726) );
  AOI22X1 U816 ( .A0(n744), .A1(n679), .B0(n681), .B1(n745), .Y(n140) );
  XNOR2X1 U817 ( .A(b[15]), .B(n680), .Y(n745) );
  XNOR2X1 U818 ( .A(n680), .B(a[4]), .Y(n836) );
  XOR2X1 U819 ( .A(b[14]), .B(n650), .Y(n744) );
  OAI22X1 U820 ( .A0(n794), .A1(n784), .B0(n782), .B1(n795), .Y(n121) );
  XNOR2X1 U821 ( .A(b[11]), .B(n653), .Y(n795) );
  XNOR2X1 U822 ( .A(n671), .B(a[10]), .Y(n837) );
  XNOR2X1 U823 ( .A(b[10]), .B(n653), .Y(n794) );
  AOI22X1 U824 ( .A0(n780), .A1(n673), .B0(n675), .B1(n781), .Y(n108) );
  XNOR2X1 U825 ( .A(b[15]), .B(n674), .Y(n781) );
  XNOR2X1 U826 ( .A(n674), .B(a[8]), .Y(n838) );
  XOR2X1 U827 ( .A(b[14]), .B(n652), .Y(n780) );
endmodule

