module CHIP( 	
	clk,
    rst_n,
    in_valid,
    in_x,
    in_y,
    move_num,
    priority_num,
    out_valid,
    out_x,
    out_y,
    move_out);

input clk,rst_n;
input in_valid;
input [2:0] in_x,in_y;
input [4:0] move_num;
input [2:0] priority_num;

output out_valid;
output [2:0] out_x,out_y;
output [4:0] move_out;

wire   C_clk;
wire   C_rst_n;
wire   C_in_valid;
wire  [2:0] C_in_x,C_in_y;
wire  [4:0] C_move_num;
wire  [2:0] C_priority_num;

wire  C_out_valid;
wire  [2:0] C_out_x,C_out_y;
wire  [4:0] C_move_out;

wire BUF_clk;
CLKBUFX20 buf0(.A(C_clk),.Y(BUF_clk));

KT I_KT(
	// Input signals
	.clk(BUF_clk),
	.rst_n(C_rst_n),
	.in_valid(C_in_valid),
	.in_x(C_in_x),
	.in_y(C_in_y),
	.move_num(C_move_num),
    .priority_num(C_priority_num),
    .out_valid(C_out_valid),
    .out_x(C_out_x),
    .out_y(C_out_y),
    .move_out(C_move_out)
);

// Input Pads
PDDDGZ I_CLK(.PAD(clk), .C(C_clk));
PDDDGZ I_RESET(.PAD(rst_n), .C(C_rst_n));
PDDDGZ I_IN_VALID(.PAD(in_valid), .C(C_in_valid));
PDDDGZ I_IN_X_2(.PAD(in_x[2]), .C(C_in_x[2]));
PDDDGZ I_IN_X_1(.PAD(in_x[1]), .C(C_in_x[1]));
PDDDGZ I_IN_X_0(.PAD(in_x[0]), .C(C_in_x[0]));
PDDDGZ I_IN_Y_2(.PAD(in_y[2]), .C(C_in_y[2]));
PDDDGZ I_IN_Y_1(.PAD(in_y[1]), .C(C_in_y[1]));
PDDDGZ I_IN_Y_0(.PAD(in_y[0]), .C(C_in_y[0]));
PDDDGZ I_MOVE_NUM_4(.PAD(move_num[4]), .C(C_move_num[4]));
PDDDGZ I_MOVE_NUM_3(.PAD(move_num[3]), .C(C_move_num[3]));
PDDDGZ I_MOVE_NUM_2(.PAD(move_num[2]), .C(C_move_num[2]));
PDDDGZ I_MOVE_NUM_1(.PAD(move_num[1]), .C(C_move_num[1]));
PDDDGZ I_MOVE_NUM_0(.PAD(move_num[0]), .C(C_move_num[0]));
PDDDGZ I_PRIORITY_NUM_2(.PAD(priority_num[2]), .C(C_priority_num[2]));
PDDDGZ I_PRIORITY_NUM_1(.PAD(priority_num[1]), .C(C_priority_num[1]));
PDDDGZ I_PRIORITY_NUM_0(.PAD(priority_num[0]), .C(C_priority_num[0]));
// Output Pads
PDD08SDGZ O_OUT_VALID(.OEN(1'b0), .I(C_out_valid), .PAD(out_valid), .C());
PDD08SDGZ O_OUT_X_0(.OEN(1'b0), .I(C_out_x[0]), .PAD(out_x[0]), .C());
PDD08SDGZ O_OUT_X_1(.OEN(1'b0), .I(C_out_x[1]), .PAD(out_x[1]), .C());
PDD08SDGZ O_OUT_X_2(.OEN(1'b0), .I(C_out_x[2]), .PAD(out_x[2]), .C());
PDD08SDGZ O_OUT_Y_0(.OEN(1'b0), .I(C_out_y[0]), .PAD(out_y[0]), .C());
PDD08SDGZ O_OUT_Y_1(.OEN(1'b0), .I(C_out_y[1]), .PAD(out_y[1]), .C());
PDD08SDGZ O_OUT_Y_2(.OEN(1'b0), .I(C_out_y[2]), .PAD(out_y[2]), .C());
PDD08SDGZ O_MOVE_OUT_0(.OEN(1'b0), .I(C_move_out[0]), .PAD(move_out[0]), .C());
PDD08SDGZ O_MOVE_OUT_1(.OEN(1'b0), .I(C_move_out[1]), .PAD(move_out[1]), .C());
PDD08SDGZ O_MOVE_OUT_2(.OEN(1'b0), .I(C_move_out[2]), .PAD(move_out[2]), .C());
PDD08SDGZ O_MOVE_OUT_3(.OEN(1'b0), .I(C_move_out[3]), .PAD(move_out[3]), .C());
PDD08SDGZ O_MOVE_OUT_4(.OEN(1'b0), .I(C_move_out[4]), .PAD(move_out[4]), .C());

// IO power 
PVDD2DGZ VDDP0 ();
PVSS2DGZ GNDP0 ();
PVDD2DGZ VDDP1 ();
PVSS2DGZ GNDP1 ();
PVDD2DGZ VDDP2 ();
PVSS2DGZ GNDP2 ();
PVDD2DGZ VDDP3 ();
PVSS2DGZ GNDP3 ();


// Core power
PVDD1DGZ VDDC0 ();
PVSS1DGZ GNDC0 ();
PVDD1DGZ VDDC1 ();
PVSS1DGZ GNDC1 ();
PVDD1DGZ VDDC2 ();
PVSS1DGZ GNDC2 ();
PVDD1DGZ VDDC3 ();
PVSS1DGZ GNDC3 ();


endmodule
/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : O-2018.06-SP1
// Date      : Mon Oct 28 10:39:52 2024
/////////////////////////////////////////////////////////////


module KT ( clk, rst_n, in_valid, in_x, in_y, move_num, priority_num, 
        out_valid, out_x, out_y, move_out );
  input [2:0] in_x;
  input [2:0] in_y;
  input [4:0] move_num;
  input [2:0] priority_num;
  output [2:0] out_x;
  output [2:0] out_y;
  output [4:0] move_out;
  input clk, rst_n, in_valid;
  output out_valid;
  wire   N2025, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931;
  wire   [4:1] cnt;
  wire   [199:0] have_tried_direction;
  wire   [74:0] x;
  wire   [74:0] y;
  wire   [1:0] cs;
  wire   [2:0] direction;
  wire   [2:0] pri;

  DFFSX1 have_tried_direction_reg_0__0_ ( .D(n1600), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[0]) );
  DFFSX1 direction_reg_1_ ( .D(n1599), .CK(clk), .SN(rst_n), .Q(n2879), .QN(
        direction[1]) );
  DFFSX1 direction_reg_2_ ( .D(n1598), .CK(clk), .SN(rst_n), .Q(n2878), .QN(
        direction[2]) );
  DFFSX1 cs_reg_0_ ( .D(n1596), .CK(clk), .SN(rst_n), .QN(cs[0]) );
  DFFSX1 cs_reg_1_ ( .D(n1594), .CK(clk), .SN(rst_n), .Q(n2925), .QN(cs[1]) );
  DFFSX1 cnt_reg_4_ ( .D(n1593), .CK(clk), .SN(rst_n), .Q(n2862), .QN(cnt[4])
         );
  DFFSX1 pri_reg_0_ ( .D(n1589), .CK(clk), .SN(rst_n), .Q(n2924), .QN(pri[0])
         );
  DFFSX1 pri_reg_2_ ( .D(n1588), .CK(clk), .SN(rst_n), .QN(pri[2]) );
  DFFSX1 pri_reg_1_ ( .D(n1587), .CK(clk), .SN(rst_n), .QN(pri[1]) );
  DFFSX1 direction_reg_0_ ( .D(n1585), .CK(clk), .SN(rst_n), .Q(n2864), .QN(
        direction[0]) );
  DFFSX1 have_tried_direction_reg_0__1_ ( .D(n1579), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[1]) );
  DFFSX1 have_tried_direction_reg_0__2_ ( .D(n1578), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[2]) );
  DFFSX1 have_tried_direction_reg_0__3_ ( .D(n1577), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[3]) );
  DFFSX1 have_tried_direction_reg_0__4_ ( .D(n1576), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[4]) );
  DFFSX1 have_tried_direction_reg_0__5_ ( .D(n1575), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[5]) );
  DFFSX1 have_tried_direction_reg_0__6_ ( .D(n1574), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[6]) );
  DFFSX1 have_tried_direction_reg_0__7_ ( .D(n1573), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[7]) );
  DFFSX1 have_tried_direction_reg_1__0_ ( .D(n1572), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[8]) );
  DFFSX1 have_tried_direction_reg_1__1_ ( .D(n1571), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[9]) );
  DFFSX1 have_tried_direction_reg_1__2_ ( .D(n1570), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[10]) );
  DFFSX1 have_tried_direction_reg_1__3_ ( .D(n1569), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[11]) );
  DFFSX1 have_tried_direction_reg_1__4_ ( .D(n1568), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[12]) );
  DFFSX1 have_tried_direction_reg_1__5_ ( .D(n1567), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[13]) );
  DFFSX1 have_tried_direction_reg_1__6_ ( .D(n1566), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[14]) );
  DFFSX1 have_tried_direction_reg_1__7_ ( .D(n1565), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[15]) );
  DFFSX1 have_tried_direction_reg_2__0_ ( .D(n1564), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[16]) );
  DFFSX1 have_tried_direction_reg_2__1_ ( .D(n1563), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[17]) );
  DFFSX1 have_tried_direction_reg_2__2_ ( .D(n1562), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[18]) );
  DFFSX1 have_tried_direction_reg_2__3_ ( .D(n1561), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[19]) );
  DFFSX1 have_tried_direction_reg_2__4_ ( .D(n1560), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[20]) );
  DFFSX1 have_tried_direction_reg_2__5_ ( .D(n1559), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[21]) );
  DFFSX1 have_tried_direction_reg_2__6_ ( .D(n1558), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[22]) );
  DFFSX1 have_tried_direction_reg_2__7_ ( .D(n1557), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[23]) );
  DFFSX1 have_tried_direction_reg_3__0_ ( .D(n1556), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[24]) );
  DFFSX1 have_tried_direction_reg_3__1_ ( .D(n1555), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[25]) );
  DFFSX1 have_tried_direction_reg_3__2_ ( .D(n1554), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[26]) );
  DFFSX1 have_tried_direction_reg_3__3_ ( .D(n1553), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[27]) );
  DFFSX1 have_tried_direction_reg_3__4_ ( .D(n1552), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[28]) );
  DFFSX1 have_tried_direction_reg_3__5_ ( .D(n1551), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[29]) );
  DFFSX1 have_tried_direction_reg_3__6_ ( .D(n1550), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[30]) );
  DFFSX1 have_tried_direction_reg_3__7_ ( .D(n1549), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[31]) );
  DFFSX1 have_tried_direction_reg_4__0_ ( .D(n1548), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[32]) );
  DFFSX1 have_tried_direction_reg_4__1_ ( .D(n1547), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[33]) );
  DFFSX1 have_tried_direction_reg_4__2_ ( .D(n1546), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[34]) );
  DFFSX1 have_tried_direction_reg_4__3_ ( .D(n1545), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[35]) );
  DFFSX1 have_tried_direction_reg_4__4_ ( .D(n1544), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[36]) );
  DFFSX1 have_tried_direction_reg_4__5_ ( .D(n1543), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[37]) );
  DFFSX1 have_tried_direction_reg_4__6_ ( .D(n1542), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[38]) );
  DFFSX1 have_tried_direction_reg_4__7_ ( .D(n1541), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[39]) );
  DFFSX1 have_tried_direction_reg_5__0_ ( .D(n1540), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[40]) );
  DFFSX1 have_tried_direction_reg_5__1_ ( .D(n1539), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[41]) );
  DFFSX1 have_tried_direction_reg_5__2_ ( .D(n1538), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[42]) );
  DFFSX1 have_tried_direction_reg_5__3_ ( .D(n1537), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[43]) );
  DFFSX1 have_tried_direction_reg_5__4_ ( .D(n1536), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[44]) );
  DFFSX1 have_tried_direction_reg_5__5_ ( .D(n1535), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[45]) );
  DFFSX1 have_tried_direction_reg_5__6_ ( .D(n1534), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[46]) );
  DFFSX1 have_tried_direction_reg_5__7_ ( .D(n1533), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[47]) );
  DFFSX1 have_tried_direction_reg_6__0_ ( .D(n1532), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[48]) );
  DFFSX1 have_tried_direction_reg_6__1_ ( .D(n1531), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[49]) );
  DFFSX1 have_tried_direction_reg_6__2_ ( .D(n1530), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[50]) );
  DFFSX1 have_tried_direction_reg_6__3_ ( .D(n1529), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[51]) );
  DFFSX1 have_tried_direction_reg_6__4_ ( .D(n1528), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[52]) );
  DFFSX1 have_tried_direction_reg_6__5_ ( .D(n1527), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[53]) );
  DFFSX1 have_tried_direction_reg_6__6_ ( .D(n1526), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[54]) );
  DFFSX1 have_tried_direction_reg_6__7_ ( .D(n1525), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[55]) );
  DFFSX1 have_tried_direction_reg_7__0_ ( .D(n1524), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[56]) );
  DFFSX1 have_tried_direction_reg_7__1_ ( .D(n1523), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[57]) );
  DFFSX1 have_tried_direction_reg_7__2_ ( .D(n1522), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[58]) );
  DFFSX1 have_tried_direction_reg_7__3_ ( .D(n1521), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[59]) );
  DFFSX1 have_tried_direction_reg_7__4_ ( .D(n1520), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[60]) );
  DFFSX1 have_tried_direction_reg_7__5_ ( .D(n1519), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[61]) );
  DFFSX1 have_tried_direction_reg_7__6_ ( .D(n1518), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[62]) );
  DFFSX1 have_tried_direction_reg_7__7_ ( .D(n1517), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[63]) );
  DFFSX1 have_tried_direction_reg_8__0_ ( .D(n1516), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[64]) );
  DFFSX1 have_tried_direction_reg_8__1_ ( .D(n1515), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[65]) );
  DFFSX1 have_tried_direction_reg_8__2_ ( .D(n1514), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[66]) );
  DFFSX1 have_tried_direction_reg_8__3_ ( .D(n1513), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[67]) );
  DFFSX1 have_tried_direction_reg_8__4_ ( .D(n1512), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[68]) );
  DFFSX1 have_tried_direction_reg_8__5_ ( .D(n1511), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[69]) );
  DFFSX1 have_tried_direction_reg_8__6_ ( .D(n1510), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[70]) );
  DFFSX1 have_tried_direction_reg_8__7_ ( .D(n1509), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[71]) );
  DFFSX1 have_tried_direction_reg_9__0_ ( .D(n1508), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[72]) );
  DFFSX1 have_tried_direction_reg_9__1_ ( .D(n1507), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[73]) );
  DFFSX1 have_tried_direction_reg_9__2_ ( .D(n1506), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[74]) );
  DFFSX1 have_tried_direction_reg_9__3_ ( .D(n1505), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[75]) );
  DFFSX1 have_tried_direction_reg_9__4_ ( .D(n1504), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[76]) );
  DFFSX1 have_tried_direction_reg_9__5_ ( .D(n1503), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[77]) );
  DFFSX1 have_tried_direction_reg_9__6_ ( .D(n1502), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[78]) );
  DFFSX1 have_tried_direction_reg_9__7_ ( .D(n1501), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[79]) );
  DFFSX1 have_tried_direction_reg_10__0_ ( .D(n1500), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[80]) );
  DFFSX1 have_tried_direction_reg_10__1_ ( .D(n1499), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[81]) );
  DFFSX1 have_tried_direction_reg_10__2_ ( .D(n1498), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[82]) );
  DFFSX1 have_tried_direction_reg_10__3_ ( .D(n1497), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[83]) );
  DFFSX1 have_tried_direction_reg_10__4_ ( .D(n1496), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[84]) );
  DFFSX1 have_tried_direction_reg_10__5_ ( .D(n1495), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[85]) );
  DFFSX1 have_tried_direction_reg_10__6_ ( .D(n1494), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[86]) );
  DFFSX1 have_tried_direction_reg_10__7_ ( .D(n1493), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[87]) );
  DFFSX1 have_tried_direction_reg_11__0_ ( .D(n1492), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[88]) );
  DFFSX1 have_tried_direction_reg_11__1_ ( .D(n1491), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[89]) );
  DFFSX1 have_tried_direction_reg_11__2_ ( .D(n1490), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[90]) );
  DFFSX1 have_tried_direction_reg_11__3_ ( .D(n1489), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[91]) );
  DFFSX1 have_tried_direction_reg_11__4_ ( .D(n1488), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[92]) );
  DFFSX1 have_tried_direction_reg_11__5_ ( .D(n1487), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[93]) );
  DFFSX1 have_tried_direction_reg_11__6_ ( .D(n1486), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[94]) );
  DFFSX1 have_tried_direction_reg_11__7_ ( .D(n1485), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[95]) );
  DFFSX1 have_tried_direction_reg_12__0_ ( .D(n1484), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[96]) );
  DFFSX1 have_tried_direction_reg_12__1_ ( .D(n1483), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[97]) );
  DFFSX1 have_tried_direction_reg_12__2_ ( .D(n1482), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[98]) );
  DFFSX1 have_tried_direction_reg_12__3_ ( .D(n1481), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[99]) );
  DFFSX1 have_tried_direction_reg_12__4_ ( .D(n1480), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[100]) );
  DFFSX1 have_tried_direction_reg_12__5_ ( .D(n1479), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[101]) );
  DFFSX1 have_tried_direction_reg_12__6_ ( .D(n1478), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[102]) );
  DFFSX1 have_tried_direction_reg_12__7_ ( .D(n1477), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[103]) );
  DFFSX1 have_tried_direction_reg_13__0_ ( .D(n1476), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[104]) );
  DFFSX1 have_tried_direction_reg_13__1_ ( .D(n1475), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[105]) );
  DFFSX1 have_tried_direction_reg_13__2_ ( .D(n1474), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[106]) );
  DFFSX1 have_tried_direction_reg_13__3_ ( .D(n1473), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[107]) );
  DFFSX1 have_tried_direction_reg_13__4_ ( .D(n1472), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[108]) );
  DFFSX1 have_tried_direction_reg_13__5_ ( .D(n1471), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[109]) );
  DFFSX1 have_tried_direction_reg_13__6_ ( .D(n1470), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[110]) );
  DFFSX1 have_tried_direction_reg_13__7_ ( .D(n1469), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[111]) );
  DFFSX1 have_tried_direction_reg_14__0_ ( .D(n1468), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[112]) );
  DFFSX1 have_tried_direction_reg_14__1_ ( .D(n1467), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[113]) );
  DFFSX1 have_tried_direction_reg_14__2_ ( .D(n1466), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[114]) );
  DFFSX1 have_tried_direction_reg_14__3_ ( .D(n1465), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[115]) );
  DFFSX1 have_tried_direction_reg_14__4_ ( .D(n1464), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[116]) );
  DFFSX1 have_tried_direction_reg_14__5_ ( .D(n1463), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[117]) );
  DFFSX1 have_tried_direction_reg_14__6_ ( .D(n1462), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[118]) );
  DFFSX1 have_tried_direction_reg_14__7_ ( .D(n1461), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[119]) );
  DFFSX1 have_tried_direction_reg_15__0_ ( .D(n1460), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[120]) );
  DFFSX1 have_tried_direction_reg_15__1_ ( .D(n1459), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[121]) );
  DFFSX1 have_tried_direction_reg_15__2_ ( .D(n1458), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[122]) );
  DFFSX1 have_tried_direction_reg_15__3_ ( .D(n1457), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[123]) );
  DFFSX1 have_tried_direction_reg_15__4_ ( .D(n1456), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[124]) );
  DFFSX1 have_tried_direction_reg_15__5_ ( .D(n1455), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[125]) );
  DFFSX1 have_tried_direction_reg_15__6_ ( .D(n1454), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[126]) );
  DFFSX1 have_tried_direction_reg_15__7_ ( .D(n1453), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[127]) );
  DFFSX1 have_tried_direction_reg_16__0_ ( .D(n1452), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[128]) );
  DFFSX1 have_tried_direction_reg_16__1_ ( .D(n1451), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[129]) );
  DFFSX1 have_tried_direction_reg_16__2_ ( .D(n1450), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[130]) );
  DFFSX1 have_tried_direction_reg_16__3_ ( .D(n1449), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[131]) );
  DFFSX1 have_tried_direction_reg_16__4_ ( .D(n1448), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[132]) );
  DFFSX1 have_tried_direction_reg_16__5_ ( .D(n1447), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[133]) );
  DFFSX1 have_tried_direction_reg_16__6_ ( .D(n1446), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[134]) );
  DFFSX1 have_tried_direction_reg_16__7_ ( .D(n1445), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[135]) );
  DFFSX1 have_tried_direction_reg_17__0_ ( .D(n1444), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[136]) );
  DFFSX1 have_tried_direction_reg_17__1_ ( .D(n1443), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[137]) );
  DFFSX1 have_tried_direction_reg_17__2_ ( .D(n1442), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[138]) );
  DFFSX1 have_tried_direction_reg_17__3_ ( .D(n1441), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[139]) );
  DFFSX1 have_tried_direction_reg_17__4_ ( .D(n1440), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[140]) );
  DFFSX1 have_tried_direction_reg_17__5_ ( .D(n1439), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[141]) );
  DFFSX1 have_tried_direction_reg_17__6_ ( .D(n1438), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[142]) );
  DFFSX1 have_tried_direction_reg_17__7_ ( .D(n1437), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[143]) );
  DFFSX1 have_tried_direction_reg_18__0_ ( .D(n1436), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[144]) );
  DFFSX1 have_tried_direction_reg_18__1_ ( .D(n1435), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[145]) );
  DFFSX1 have_tried_direction_reg_18__2_ ( .D(n1434), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[146]) );
  DFFSX1 have_tried_direction_reg_18__3_ ( .D(n1433), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[147]) );
  DFFSX1 have_tried_direction_reg_18__4_ ( .D(n1432), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[148]) );
  DFFSX1 have_tried_direction_reg_18__5_ ( .D(n1431), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[149]) );
  DFFSX1 have_tried_direction_reg_18__6_ ( .D(n1430), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[150]) );
  DFFSX1 have_tried_direction_reg_18__7_ ( .D(n1429), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[151]) );
  DFFSX1 have_tried_direction_reg_19__0_ ( .D(n1428), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[152]) );
  DFFSX1 have_tried_direction_reg_19__1_ ( .D(n1427), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[153]) );
  DFFSX1 have_tried_direction_reg_19__2_ ( .D(n1426), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[154]) );
  DFFSX1 have_tried_direction_reg_19__3_ ( .D(n1425), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[155]) );
  DFFSX1 have_tried_direction_reg_19__4_ ( .D(n1424), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[156]) );
  DFFSX1 have_tried_direction_reg_19__5_ ( .D(n1423), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[157]) );
  DFFSX1 have_tried_direction_reg_19__6_ ( .D(n1422), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[158]) );
  DFFSX1 have_tried_direction_reg_19__7_ ( .D(n1421), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[159]) );
  DFFSX1 have_tried_direction_reg_20__0_ ( .D(n1420), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[160]) );
  DFFSX1 have_tried_direction_reg_20__1_ ( .D(n1419), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[161]) );
  DFFSX1 have_tried_direction_reg_20__2_ ( .D(n1418), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[162]) );
  DFFSX1 have_tried_direction_reg_20__3_ ( .D(n1417), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[163]) );
  DFFSX1 have_tried_direction_reg_20__4_ ( .D(n1416), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[164]) );
  DFFSX1 have_tried_direction_reg_20__5_ ( .D(n1415), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[165]) );
  DFFSX1 have_tried_direction_reg_20__6_ ( .D(n1414), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[166]) );
  DFFSX1 have_tried_direction_reg_20__7_ ( .D(n1413), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[167]) );
  DFFSX1 have_tried_direction_reg_21__0_ ( .D(n1412), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[168]) );
  DFFSX1 have_tried_direction_reg_21__1_ ( .D(n1411), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[169]) );
  DFFSX1 have_tried_direction_reg_21__2_ ( .D(n1410), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[170]) );
  DFFSX1 have_tried_direction_reg_21__3_ ( .D(n1409), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[171]) );
  DFFSX1 have_tried_direction_reg_21__4_ ( .D(n1408), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[172]) );
  DFFSX1 have_tried_direction_reg_21__5_ ( .D(n1407), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[173]) );
  DFFSX1 have_tried_direction_reg_21__6_ ( .D(n1406), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[174]) );
  DFFSX1 have_tried_direction_reg_21__7_ ( .D(n1405), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[175]) );
  DFFSX1 have_tried_direction_reg_22__0_ ( .D(n1404), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[176]) );
  DFFSX1 have_tried_direction_reg_22__1_ ( .D(n1403), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[177]) );
  DFFSX1 have_tried_direction_reg_22__2_ ( .D(n1402), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[178]) );
  DFFSX1 have_tried_direction_reg_22__3_ ( .D(n1401), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[179]) );
  DFFSX1 have_tried_direction_reg_22__4_ ( .D(n1400), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[180]) );
  DFFSX1 have_tried_direction_reg_22__5_ ( .D(n1399), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[181]) );
  DFFSX1 have_tried_direction_reg_22__6_ ( .D(n1398), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[182]) );
  DFFSX1 have_tried_direction_reg_22__7_ ( .D(n1397), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[183]) );
  DFFSX1 have_tried_direction_reg_23__0_ ( .D(n1396), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[184]) );
  DFFSX1 have_tried_direction_reg_23__1_ ( .D(n1395), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[185]) );
  DFFSX1 have_tried_direction_reg_23__2_ ( .D(n1394), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[186]) );
  DFFSX1 have_tried_direction_reg_23__3_ ( .D(n1393), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[187]) );
  DFFSX1 have_tried_direction_reg_23__4_ ( .D(n1392), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[188]) );
  DFFSX1 have_tried_direction_reg_23__5_ ( .D(n1391), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[189]) );
  DFFSX1 have_tried_direction_reg_23__6_ ( .D(n1390), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[190]) );
  DFFSX1 have_tried_direction_reg_23__7_ ( .D(n1389), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[191]) );
  DFFSX1 have_tried_direction_reg_24__0_ ( .D(n1388), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[192]) );
  DFFSX1 have_tried_direction_reg_24__1_ ( .D(n1387), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[193]) );
  DFFSX1 have_tried_direction_reg_24__2_ ( .D(n1386), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[194]) );
  DFFSX1 have_tried_direction_reg_24__3_ ( .D(n1385), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[195]) );
  DFFSX1 have_tried_direction_reg_24__4_ ( .D(n1384), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[196]) );
  DFFSX1 have_tried_direction_reg_24__5_ ( .D(n1383), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[197]) );
  DFFSX1 have_tried_direction_reg_24__6_ ( .D(n1382), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[198]) );
  DFFSX1 have_tried_direction_reg_24__7_ ( .D(n1381), .CK(clk), .SN(rst_n), 
        .QN(have_tried_direction[199]) );
  DFFSX1 y_reg_0__2_ ( .D(n1752), .CK(clk), .SN(rst_n), .Q(y[2]), .QN(n2913)
         );
  DFFSX1 y_reg_1__2_ ( .D(n1749), .CK(clk), .SN(rst_n), .Q(y[5]), .QN(n2912)
         );
  DFFSX1 y_reg_2__2_ ( .D(n1746), .CK(clk), .SN(rst_n), .Q(y[8]), .QN(n2923)
         );
  DFFSX1 y_reg_3__2_ ( .D(n1743), .CK(clk), .SN(rst_n), .Q(y[11]), .QN(n2906)
         );
  DFFSX1 y_reg_4__2_ ( .D(n1740), .CK(clk), .SN(rst_n), .Q(y[14]), .QN(n2918)
         );
  DFFSX1 y_reg_5__2_ ( .D(n1737), .CK(clk), .SN(rst_n), .Q(y[17]), .QN(n2869)
         );
  DFFSX1 y_reg_6__2_ ( .D(n1734), .CK(clk), .SN(rst_n), .Q(y[20]), .QN(n2919)
         );
  DFFSX1 y_reg_7__2_ ( .D(n1731), .CK(clk), .SN(rst_n), .Q(y[23]), .QN(n2866)
         );
  DFFSX1 y_reg_8__2_ ( .D(n1728), .CK(clk), .SN(rst_n), .Q(y[26]), .QN(n2916)
         );
  DFFSX1 y_reg_9__2_ ( .D(n1725), .CK(clk), .SN(rst_n), .Q(y[29]), .QN(n2917)
         );
  DFFSX1 y_reg_10__2_ ( .D(n1722), .CK(clk), .SN(rst_n), .Q(y[32]), .QN(n2868)
         );
  DFFSX1 y_reg_11__2_ ( .D(n1719), .CK(clk), .SN(rst_n), .Q(y[35]), .QN(n2870)
         );
  DFFSX1 y_reg_12__2_ ( .D(n1716), .CK(clk), .SN(rst_n), .Q(y[38]), .QN(n2920)
         );
  DFFSX1 y_reg_13__2_ ( .D(n1713), .CK(clk), .SN(rst_n), .Q(y[41]), .QN(n2871)
         );
  DFFSX1 y_reg_14__2_ ( .D(n1710), .CK(clk), .SN(rst_n), .Q(y[44]), .QN(n2921)
         );
  DFFSX1 y_reg_15__2_ ( .D(n1707), .CK(clk), .SN(rst_n), .Q(y[47]), .QN(n2914)
         );
  DFFSX1 y_reg_16__2_ ( .D(n1704), .CK(clk), .SN(rst_n), .Q(y[50]), .QN(n2865)
         );
  DFFSX1 y_reg_17__2_ ( .D(n1701), .CK(clk), .SN(rst_n), .Q(y[53]), .QN(n2867)
         );
  DFFSX1 y_reg_18__2_ ( .D(n1698), .CK(clk), .SN(rst_n), .Q(y[56]), .QN(n2907)
         );
  DFFSX1 y_reg_19__2_ ( .D(n1695), .CK(clk), .SN(rst_n), .Q(y[59]), .QN(n2909)
         );
  DFFSX1 y_reg_20__2_ ( .D(n1692), .CK(clk), .SN(rst_n), .Q(y[62]), .QN(n2922)
         );
  DFFSX1 y_reg_21__2_ ( .D(n1689), .CK(clk), .SN(rst_n), .Q(y[65]), .QN(n2872)
         );
  DFFSX1 y_reg_22__2_ ( .D(n1686), .CK(clk), .SN(rst_n), .Q(y[68]), .QN(n2915)
         );
  DFFSX1 y_reg_23__2_ ( .D(n1683), .CK(clk), .SN(rst_n), .Q(y[71]) );
  DFFSX1 y_reg_24__2_ ( .D(n1680), .CK(clk), .SN(rst_n), .Q(y[74]), .QN(n2908)
         );
  DFFSX1 x_reg_0__0_ ( .D(n1679), .CK(clk), .SN(rst_n), .Q(x[0]) );
  DFFSX1 x_reg_1__0_ ( .D(n1676), .CK(clk), .SN(rst_n), .Q(x[3]) );
  DFFSX1 x_reg_2__0_ ( .D(n1673), .CK(clk), .SN(rst_n), .Q(x[6]) );
  DFFSX1 x_reg_3__0_ ( .D(n1670), .CK(clk), .SN(rst_n), .Q(x[9]), .QN(n2929)
         );
  DFFSX1 x_reg_4__0_ ( .D(n1667), .CK(clk), .SN(rst_n), .Q(x[12]) );
  DFFSX1 x_reg_5__0_ ( .D(n1664), .CK(clk), .SN(rst_n), .Q(x[15]) );
  DFFSX1 x_reg_6__0_ ( .D(n1661), .CK(clk), .SN(rst_n), .Q(x[18]) );
  DFFSX1 x_reg_7__0_ ( .D(n1658), .CK(clk), .SN(rst_n), .Q(x[21]) );
  DFFSX1 x_reg_8__0_ ( .D(n1655), .CK(clk), .SN(rst_n), .Q(x[24]) );
  DFFSX1 x_reg_9__0_ ( .D(n1652), .CK(clk), .SN(rst_n), .Q(x[27]) );
  DFFSX1 x_reg_10__0_ ( .D(n1649), .CK(clk), .SN(rst_n), .Q(x[30]) );
  DFFSX1 x_reg_11__0_ ( .D(n1646), .CK(clk), .SN(rst_n), .Q(x[33]) );
  DFFSX1 x_reg_12__0_ ( .D(n1643), .CK(clk), .SN(rst_n), .Q(x[36]) );
  DFFSX1 x_reg_13__0_ ( .D(n1640), .CK(clk), .SN(rst_n), .Q(x[39]) );
  DFFSX1 x_reg_14__0_ ( .D(n1637), .CK(clk), .SN(rst_n), .Q(x[42]) );
  DFFSX1 x_reg_15__0_ ( .D(n1634), .CK(clk), .SN(rst_n), .Q(x[45]) );
  DFFSX1 x_reg_16__0_ ( .D(n1631), .CK(clk), .SN(rst_n), .Q(x[48]) );
  DFFSX1 x_reg_17__0_ ( .D(n1628), .CK(clk), .SN(rst_n), .Q(x[51]) );
  DFFSX1 x_reg_18__0_ ( .D(n1625), .CK(clk), .SN(rst_n), .Q(x[54]) );
  DFFSX1 x_reg_19__0_ ( .D(n1622), .CK(clk), .SN(rst_n), .Q(x[57]) );
  DFFSX1 x_reg_20__0_ ( .D(n1619), .CK(clk), .SN(rst_n), .Q(x[60]) );
  DFFSX1 x_reg_21__0_ ( .D(n1616), .CK(clk), .SN(rst_n), .Q(x[63]) );
  DFFSX1 x_reg_22__0_ ( .D(n1613), .CK(clk), .SN(rst_n), .Q(x[66]) );
  DFFSX1 x_reg_23__0_ ( .D(n1610), .CK(clk), .SN(rst_n), .Q(x[69]), .QN(n2905)
         );
  DFFSX1 x_reg_24__0_ ( .D(n1607), .CK(clk), .SN(rst_n), .Q(x[72]), .QN(n2911)
         );
  DFFSX1 y_reg_0__0_ ( .D(n1754), .CK(clk), .SN(rst_n), .Q(y[0]), .QN(n2883)
         );
  DFFSX1 y_reg_1__0_ ( .D(n1751), .CK(clk), .SN(rst_n), .Q(y[3]), .QN(n2894)
         );
  DFFSX1 y_reg_2__0_ ( .D(n1748), .CK(clk), .SN(rst_n), .Q(y[6]), .QN(n2897)
         );
  DFFSX1 y_reg_3__0_ ( .D(n1745), .CK(clk), .SN(rst_n), .Q(y[9]), .QN(n2881)
         );
  DFFSX1 y_reg_4__0_ ( .D(n1742), .CK(clk), .SN(rst_n), .Q(y[12]), .QN(n2898)
         );
  DFFSX1 y_reg_5__0_ ( .D(n1739), .CK(clk), .SN(rst_n), .Q(y[15]), .QN(n2890)
         );
  DFFSX1 y_reg_6__0_ ( .D(n1736), .CK(clk), .SN(rst_n), .Q(y[18]), .QN(n2899)
         );
  DFFSX1 y_reg_7__0_ ( .D(n1733), .CK(clk), .SN(rst_n), .Q(y[21]), .QN(n2884)
         );
  DFFSX1 y_reg_8__0_ ( .D(n1730), .CK(clk), .SN(rst_n), .Q(y[24]), .QN(n2889)
         );
  DFFSX1 y_reg_9__0_ ( .D(n1727), .CK(clk), .SN(rst_n), .Q(y[27]), .QN(n2896)
         );
  DFFSX1 y_reg_10__0_ ( .D(n1724), .CK(clk), .SN(rst_n), .Q(y[30]), .QN(n2900)
         );
  DFFSX1 y_reg_11__0_ ( .D(n1721), .CK(clk), .SN(rst_n), .Q(y[33]), .QN(n2891)
         );
  DFFSX1 y_reg_12__0_ ( .D(n1718), .CK(clk), .SN(rst_n), .Q(y[36]), .QN(n2901)
         );
  DFFSX1 y_reg_13__0_ ( .D(n1715), .CK(clk), .SN(rst_n), .Q(y[39]), .QN(n2892)
         );
  DFFSX1 y_reg_14__0_ ( .D(n1712), .CK(clk), .SN(rst_n), .Q(y[42]), .QN(n2902)
         );
  DFFSX1 y_reg_15__0_ ( .D(n1709), .CK(clk), .SN(rst_n), .Q(y[45]), .QN(n2885)
         );
  DFFSX1 y_reg_16__0_ ( .D(n1706), .CK(clk), .SN(rst_n), .Q(y[48]), .QN(n2882)
         );
  DFFSX1 y_reg_17__0_ ( .D(n1703), .CK(clk), .SN(rst_n), .Q(y[51]), .QN(n2888)
         );
  DFFSX1 y_reg_18__0_ ( .D(n1700), .CK(clk), .SN(rst_n), .Q(y[54]), .QN(n2903)
         );
  DFFSX1 y_reg_19__0_ ( .D(n1697), .CK(clk), .SN(rst_n), .Q(y[57]), .QN(n2893)
         );
  DFFSX1 y_reg_20__0_ ( .D(n1694), .CK(clk), .SN(rst_n), .Q(y[60]), .QN(n2904)
         );
  DFFSX1 y_reg_21__0_ ( .D(n1691), .CK(clk), .SN(rst_n), .Q(y[63]), .QN(n2887)
         );
  DFFSX1 y_reg_22__0_ ( .D(n1688), .CK(clk), .SN(rst_n), .Q(y[66]), .QN(n2895)
         );
  DFFSX1 y_reg_23__0_ ( .D(n1685), .CK(clk), .SN(rst_n), .Q(y[69]) );
  DFFSX1 y_reg_24__0_ ( .D(n1682), .CK(clk), .SN(rst_n), .Q(y[72]), .QN(n2886)
         );
  DFFSX1 y_reg_0__1_ ( .D(n1753), .CK(clk), .SN(rst_n), .Q(y[1]) );
  DFFSX1 y_reg_1__1_ ( .D(n1750), .CK(clk), .SN(rst_n), .Q(y[4]) );
  DFFSX1 y_reg_2__1_ ( .D(n1747), .CK(clk), .SN(rst_n), .Q(y[7]) );
  DFFSX1 y_reg_3__1_ ( .D(n1744), .CK(clk), .SN(rst_n), .Q(y[10]), .QN(n2928)
         );
  DFFSX1 y_reg_4__1_ ( .D(n1741), .CK(clk), .SN(rst_n), .Q(y[13]) );
  DFFSX1 y_reg_5__1_ ( .D(n1738), .CK(clk), .SN(rst_n), .Q(y[16]) );
  DFFSX1 y_reg_6__1_ ( .D(n1735), .CK(clk), .SN(rst_n), .Q(y[19]) );
  DFFSX1 y_reg_7__1_ ( .D(n1732), .CK(clk), .SN(rst_n), .Q(y[22]) );
  DFFSX1 y_reg_8__1_ ( .D(n1729), .CK(clk), .SN(rst_n), .Q(y[25]) );
  DFFSX1 y_reg_9__1_ ( .D(n1726), .CK(clk), .SN(rst_n), .Q(y[28]) );
  DFFSX1 y_reg_10__1_ ( .D(n1723), .CK(clk), .SN(rst_n), .Q(y[31]) );
  DFFSX1 y_reg_11__1_ ( .D(n1720), .CK(clk), .SN(rst_n), .Q(y[34]) );
  DFFSX1 y_reg_12__1_ ( .D(n1717), .CK(clk), .SN(rst_n), .Q(y[37]) );
  DFFSX1 y_reg_13__1_ ( .D(n1714), .CK(clk), .SN(rst_n), .Q(y[40]) );
  DFFSX1 y_reg_14__1_ ( .D(n1711), .CK(clk), .SN(rst_n), .Q(y[43]) );
  DFFSX1 y_reg_15__1_ ( .D(n1708), .CK(clk), .SN(rst_n), .Q(y[46]) );
  DFFSX1 y_reg_16__1_ ( .D(n1705), .CK(clk), .SN(rst_n), .Q(y[49]) );
  DFFSX1 y_reg_17__1_ ( .D(n1702), .CK(clk), .SN(rst_n), .Q(y[52]) );
  DFFSX1 y_reg_18__1_ ( .D(n1699), .CK(clk), .SN(rst_n), .Q(y[55]) );
  DFFSX1 y_reg_19__1_ ( .D(n1696), .CK(clk), .SN(rst_n), .Q(y[58]) );
  DFFSX1 y_reg_20__1_ ( .D(n1693), .CK(clk), .SN(rst_n), .Q(y[61]) );
  DFFSX1 y_reg_21__1_ ( .D(n1690), .CK(clk), .SN(rst_n), .Q(y[64]) );
  DFFSX1 y_reg_22__1_ ( .D(n1687), .CK(clk), .SN(rst_n), .Q(y[67]) );
  DFFSX1 y_reg_23__1_ ( .D(n1684), .CK(clk), .SN(rst_n), .Q(y[70]) );
  DFFSX1 y_reg_24__1_ ( .D(n1681), .CK(clk), .SN(rst_n), .Q(y[73]), .QN(n2910)
         );
  DFFSX1 x_reg_0__1_ ( .D(n1678), .CK(clk), .SN(rst_n), .Q(x[1]) );
  DFFSX1 x_reg_1__1_ ( .D(n1675), .CK(clk), .SN(rst_n), .Q(x[4]) );
  DFFSX1 x_reg_2__1_ ( .D(n1672), .CK(clk), .SN(rst_n), .Q(x[7]) );
  DFFSX1 x_reg_3__1_ ( .D(n1669), .CK(clk), .SN(rst_n), .Q(x[10]), .QN(n2931)
         );
  DFFSX1 x_reg_4__1_ ( .D(n1666), .CK(clk), .SN(rst_n), .Q(x[13]) );
  DFFSX1 x_reg_5__1_ ( .D(n1663), .CK(clk), .SN(rst_n), .Q(x[16]) );
  DFFSX1 x_reg_6__1_ ( .D(n1660), .CK(clk), .SN(rst_n), .Q(x[19]) );
  DFFSX1 x_reg_7__1_ ( .D(n1657), .CK(clk), .SN(rst_n), .Q(x[22]) );
  DFFSX1 x_reg_8__1_ ( .D(n1654), .CK(clk), .SN(rst_n), .Q(x[25]) );
  DFFSX1 x_reg_9__1_ ( .D(n1651), .CK(clk), .SN(rst_n), .Q(x[28]) );
  DFFSX1 x_reg_10__1_ ( .D(n1648), .CK(clk), .SN(rst_n), .Q(x[31]) );
  DFFSX1 x_reg_11__1_ ( .D(n1645), .CK(clk), .SN(rst_n), .Q(x[34]) );
  DFFSX1 x_reg_12__1_ ( .D(n1642), .CK(clk), .SN(rst_n), .Q(x[37]) );
  DFFSX1 x_reg_13__1_ ( .D(n1639), .CK(clk), .SN(rst_n), .Q(x[40]) );
  DFFSX1 x_reg_14__1_ ( .D(n1636), .CK(clk), .SN(rst_n), .Q(x[43]) );
  DFFSX1 x_reg_15__1_ ( .D(n1633), .CK(clk), .SN(rst_n), .Q(x[46]) );
  DFFSX1 x_reg_16__1_ ( .D(n1630), .CK(clk), .SN(rst_n), .Q(x[49]) );
  DFFSX1 x_reg_17__1_ ( .D(n1627), .CK(clk), .SN(rst_n), .Q(x[52]) );
  DFFSX1 x_reg_18__1_ ( .D(n1624), .CK(clk), .SN(rst_n), .Q(x[55]) );
  DFFSX1 x_reg_19__1_ ( .D(n1621), .CK(clk), .SN(rst_n), .Q(x[58]) );
  DFFSX1 x_reg_20__1_ ( .D(n1618), .CK(clk), .SN(rst_n), .Q(x[61]) );
  DFFSX1 x_reg_21__1_ ( .D(n1615), .CK(clk), .SN(rst_n), .Q(x[64]) );
  DFFSX1 x_reg_22__1_ ( .D(n1612), .CK(clk), .SN(rst_n), .Q(x[67]) );
  DFFSX1 x_reg_23__1_ ( .D(n1609), .CK(clk), .SN(rst_n), .Q(x[70]) );
  DFFSX1 x_reg_24__1_ ( .D(n1606), .CK(clk), .SN(rst_n), .Q(x[73]), .QN(n2877)
         );
  DFFSX1 x_reg_24__2_ ( .D(n1755), .CK(clk), .SN(rst_n), .Q(x[74]), .QN(n2880)
         );
  DFFSX1 x_reg_0__2_ ( .D(n1677), .CK(clk), .SN(rst_n), .Q(x[2]) );
  DFFSX1 x_reg_1__2_ ( .D(n1674), .CK(clk), .SN(rst_n), .Q(x[5]) );
  DFFSX1 x_reg_2__2_ ( .D(n1671), .CK(clk), .SN(rst_n), .Q(x[8]) );
  DFFSX1 x_reg_3__2_ ( .D(n1668), .CK(clk), .SN(rst_n), .Q(x[11]), .QN(n2930)
         );
  DFFSX1 x_reg_4__2_ ( .D(n1665), .CK(clk), .SN(rst_n), .Q(x[14]) );
  DFFSX1 x_reg_5__2_ ( .D(n1662), .CK(clk), .SN(rst_n), .Q(x[17]) );
  DFFSX1 x_reg_6__2_ ( .D(n1659), .CK(clk), .SN(rst_n), .Q(x[20]) );
  DFFSX1 x_reg_7__2_ ( .D(n1656), .CK(clk), .SN(rst_n), .Q(x[23]) );
  DFFSX1 x_reg_8__2_ ( .D(n1653), .CK(clk), .SN(rst_n), .Q(x[26]) );
  DFFSX1 x_reg_9__2_ ( .D(n1650), .CK(clk), .SN(rst_n), .Q(x[29]) );
  DFFSX1 x_reg_10__2_ ( .D(n1647), .CK(clk), .SN(rst_n), .Q(x[32]) );
  DFFSX1 x_reg_11__2_ ( .D(n1644), .CK(clk), .SN(rst_n), .Q(x[35]) );
  DFFSX1 x_reg_12__2_ ( .D(n1641), .CK(clk), .SN(rst_n), .Q(x[38]) );
  DFFSX1 x_reg_13__2_ ( .D(n1638), .CK(clk), .SN(rst_n), .Q(x[41]) );
  DFFSX1 x_reg_14__2_ ( .D(n1635), .CK(clk), .SN(rst_n), .Q(x[44]) );
  DFFSX1 x_reg_15__2_ ( .D(n1632), .CK(clk), .SN(rst_n), .Q(x[47]) );
  DFFSX1 x_reg_16__2_ ( .D(n1629), .CK(clk), .SN(rst_n), .Q(x[50]) );
  DFFSX1 x_reg_17__2_ ( .D(n1626), .CK(clk), .SN(rst_n), .Q(x[53]) );
  DFFSX1 x_reg_18__2_ ( .D(n1623), .CK(clk), .SN(rst_n), .Q(x[56]) );
  DFFSX1 x_reg_19__2_ ( .D(n1620), .CK(clk), .SN(rst_n), .Q(x[59]) );
  DFFSX1 x_reg_20__2_ ( .D(n1617), .CK(clk), .SN(rst_n), .Q(x[62]) );
  DFFSX1 x_reg_21__2_ ( .D(n1614), .CK(clk), .SN(rst_n), .Q(x[65]) );
  DFFSX1 x_reg_22__2_ ( .D(n1611), .CK(clk), .SN(rst_n), .Q(x[68]) );
  DFFSX1 x_reg_23__2_ ( .D(n1608), .CK(clk), .SN(rst_n), .Q(x[71]) );
  DFFSX1 cnt_out_reg_1_ ( .D(n1604), .CK(clk), .SN(rst_n), .Q(n2927), .QN(
        move_out[1]) );
  DFFSX1 cnt_out_reg_4_ ( .D(n1601), .CK(clk), .SN(rst_n), .Q(n2926), .QN(
        move_out[4]) );
  DFFSX1 cnt_out_reg_0_ ( .D(n1605), .CK(clk), .SN(rst_n), .Q(n2874), .QN(
        move_out[0]) );
  DFFSX1 cnt_out_reg_3_ ( .D(n1602), .CK(clk), .SN(rst_n), .Q(n2873), .QN(
        move_out[3]) );
  DFFSX1 cnt_reg_0_ ( .D(n1592), .CK(clk), .SN(rst_n), .Q(n2863), .QN(N2025)
         );
  DFFSX1 out_valid_reg ( .D(n1595), .CK(clk), .SN(rst_n), .QN(out_valid) );
  DFFSX1 out_y_reg_2_ ( .D(n1586), .CK(clk), .SN(rst_n), .QN(out_y[2]) );
  DFFSX1 out_x_reg_0_ ( .D(n1584), .CK(clk), .SN(rst_n), .QN(out_x[0]) );
  DFFSX1 out_y_reg_0_ ( .D(n1583), .CK(clk), .SN(rst_n), .QN(out_y[0]) );
  DFFSX1 out_y_reg_1_ ( .D(n1582), .CK(clk), .SN(rst_n), .QN(out_y[1]) );
  DFFSX1 out_x_reg_1_ ( .D(n1581), .CK(clk), .SN(rst_n), .QN(out_x[1]) );
  DFFSX1 out_x_reg_2_ ( .D(n1580), .CK(clk), .SN(rst_n), .QN(out_x[2]) );
  DFFSX1 cnt_reg_2_ ( .D(n1590), .CK(clk), .SN(rst_n), .Q(n2875), .QN(cnt[2])
         );
  DFFSX1 cnt_reg_1_ ( .D(n1591), .CK(clk), .SN(rst_n), .Q(n2876), .QN(cnt[1])
         );
  DFFSX2 cnt_out_reg_2_ ( .D(n1603), .CK(clk), .SN(rst_n), .QN(move_out[2]) );
  DFFSX2 cnt_reg_3_ ( .D(n1597), .CK(clk), .SN(rst_n), .Q(n2861), .QN(cnt[3])
         );
  BUFX3 U1755 ( .A(n2852), .Y(n1769) );
  BUFX3 U1756 ( .A(n1811), .Y(n1978) );
  AOI211X2 U1757 ( .A0(cnt[4]), .A1(n2790), .B0(n2674), .C0(n2699), .Y(n2842)
         );
  BUFX3 U1758 ( .A(n1849), .Y(n1968) );
  INVX1 U1759 ( .A(n1885), .Y(n1764) );
  CLKBUFX3 U1760 ( .A(n2796), .Y(n2811) );
  CLKBUFX3 U1761 ( .A(n2687), .Y(n2692) );
  CLKBUFX3 U1762 ( .A(n2802), .Y(n2824) );
  CLKBUFX3 U1763 ( .A(n2690), .Y(n2691) );
  CLKBUFX3 U1764 ( .A(n2788), .Y(n2812) );
  CLKBUFX3 U1765 ( .A(n2677), .Y(n2813) );
  CLKINVX3 U1766 ( .A(n1769), .Y(n2638) );
  NOR2X1 U1767 ( .A(n2853), .B(n2390), .Y(n2852) );
  INVX2 U1768 ( .A(n1764), .Y(n2798) );
  INVX4 U1769 ( .A(n1764), .Y(n1757) );
  AOI221X1 U1770 ( .A0(n2524), .A1(n1884), .B0(n1883), .B1(n1882), .C0(n1881), 
        .Y(n1885) );
  INVX8 U1771 ( .A(n2219), .Y(n1758) );
  CLKINVX8 U1772 ( .A(n2685), .Y(n1759) );
  CLKINVX2 U1773 ( .A(n2634), .Y(n2703) );
  CLKINVX2 U1774 ( .A(n2631), .Y(n2761) );
  CLKINVX2 U1775 ( .A(n2637), .Y(n2711) );
  CLKINVX2 U1776 ( .A(n2629), .Y(n2707) );
  CLKINVX4 U1777 ( .A(n2776), .Y(n1765) );
  CLKBUFX3 U1778 ( .A(n2624), .Y(n2587) );
  NOR2X2 U1779 ( .A(n2862), .B(n2752), .Y(n2192) );
  CLKBUFX3 U1780 ( .A(n2623), .Y(n2583) );
  NOR2X2 U1781 ( .A(n2862), .B(n2578), .Y(n2193) );
  AOI22X1 U1782 ( .A0(n1766), .A1(n2861), .B0(cnt[3]), .B1(n2790), .Y(n2678)
         );
  CLKBUFX3 U1783 ( .A(n2622), .Y(n2577) );
  CLKINVX2 U1784 ( .A(n2640), .Y(n2684) );
  CLKBUFX3 U1785 ( .A(n2625), .Y(n2584) );
  CLKINVX8 U1786 ( .A(n2790), .Y(n1766) );
  INVX8 U1787 ( .A(n2578), .Y(n1760) );
  CLKINVX8 U1788 ( .A(n2752), .Y(n1761) );
  INVX2 U1789 ( .A(n1854), .Y(n2776) );
  INVX8 U1790 ( .A(n2735), .Y(n1762) );
  INVX8 U1791 ( .A(n2732), .Y(n1763) );
  OAI32XL U1792 ( .A0(N2025), .A1(n2720), .A2(n2838), .B0(n2849), .B1(n2863), 
        .Y(n1592) );
  AND2XL U1793 ( .A(n2755), .B(n2638), .Y(n2657) );
  CLKINVX4 U1794 ( .A(n2628), .Y(n2662) );
  AND2XL U1795 ( .A(n2743), .B(n2638), .Y(n2647) );
  AOI211XL U1796 ( .A0(n2861), .A1(n2732), .B0(n2847), .C0(n2840), .Y(n2680)
         );
  OAI221XL U1797 ( .A0(n2840), .A1(cnt[4]), .B0(n2839), .B1(n2862), .C0(n2838), 
        .Y(n2841) );
  AOI222XL U1798 ( .A0(n2864), .A1(n2854), .B0(n2853), .B1(pri[0]), .C0(n1769), 
        .C1(n2851), .Y(n2858) );
  NOR2X1 U1799 ( .A(n2268), .B(n2267), .Y(n2853) );
  NOR2XL U1800 ( .A(n2688), .B(n2054), .Y(n2055) );
  AOI2BB1XL U1801 ( .A0N(n2923), .A1N(n2216), .B0(n2215), .Y(n2226) );
  AND4XL U1802 ( .A(n2253), .B(n2252), .C(n2251), .D(n2250), .Y(n2254) );
  OR2XL U1803 ( .A(n2546), .B(n2558), .Y(n2544) );
  AND2XL U1804 ( .A(n2541), .B(n2536), .Y(n2533) );
  MXI2XL U1805 ( .A(n1873), .B(n1877), .S0(n1847), .Y(n1848) );
  NOR2X1 U1806 ( .A(n2274), .B(n2273), .Y(n2390) );
  MXI2XL U1807 ( .A(n1930), .B(n1929), .S0(n1809), .Y(n1810) );
  NOR2X1 U1808 ( .A(n2210), .B(n2209), .Y(n2274) );
  OR2XL U1809 ( .A(n1877), .B(n2521), .Y(n1871) );
  INVXL U1810 ( .A(n2521), .Y(n1878) );
  INVXL U1811 ( .A(n2512), .Y(n1872) );
  INVXL U1812 ( .A(n1916), .Y(n1867) );
  AND4XL U1813 ( .A(n2062), .B(n2061), .C(n2060), .D(n2059), .Y(n2073) );
  AND4XL U1814 ( .A(n2188), .B(n2187), .C(n2186), .D(n2185), .Y(n2202) );
  AND4XL U1815 ( .A(n2111), .B(n2110), .C(n2109), .D(n2108), .Y(n2121) );
  NOR2X1 U1816 ( .A(n2842), .B(n2678), .Y(n1916) );
  AND4XL U1817 ( .A(n2079), .B(n2078), .C(n2077), .D(n2076), .Y(n2089) );
  AND4XL U1818 ( .A(n2095), .B(n2094), .C(n2093), .D(n2092), .Y(n2105) );
  AND4XL U1819 ( .A(n2147), .B(n2146), .C(n2145), .D(n2144), .Y(n2157) );
  AND4XL U1820 ( .A(n2131), .B(n2130), .C(n2129), .D(n2128), .Y(n2141) );
  INVX1 U1821 ( .A(n2842), .Y(n1778) );
  AND4XL U1822 ( .A(n2163), .B(n2162), .C(n2161), .D(n2160), .Y(n2173) );
  AOI221XL U1823 ( .A0(direction[0]), .A1(pri[0]), .B0(n2864), .B1(n2924), 
        .C0(n2272), .Y(n2273) );
  AND2XL U1824 ( .A(priority_num[1]), .B(n2855), .Y(n2552) );
  AOI31XL U1825 ( .A0(cs[0]), .A1(n2925), .A2(n2671), .B0(n2278), .Y(n1594) );
  INVX2 U1826 ( .A(n2635), .Y(n2699) );
  INVX2 U1827 ( .A(n2727), .Y(n2738) );
  AOI31XL U1828 ( .A0(direction[0]), .A1(direction[1]), .A2(direction[2]), 
        .B0(n2590), .Y(n1929) );
  OR2XL U1829 ( .A(n2862), .B(n2776), .Y(n2178) );
  INVX2 U1830 ( .A(n2780), .Y(n1859) );
  NOR2X2 U1831 ( .A(n2790), .B(n2718), .Y(n2743) );
  NOR2X2 U1832 ( .A(n2790), .B(n2713), .Y(n2755) );
  NOR2XL U1833 ( .A(cnt[2]), .B(n2844), .Y(n2058) );
  CLKINVX4 U1834 ( .A(n2063), .Y(n1767) );
  NOR2X2 U1835 ( .A(cs[0]), .B(n2925), .Y(n2591) );
  INVXL U1836 ( .A(n2524), .Y(n1883) );
  AOI21XL U1837 ( .A0(n2512), .A1(n1871), .B0(n1870), .Y(n1884) );
  AOI21X1 U1838 ( .A0(n2714), .A1(n1846), .B0(n1845), .Y(n2521) );
  NAND4XL U1839 ( .A(n1833), .B(n1832), .C(n1831), .D(n1830), .Y(n1846) );
  OAI21XL U1840 ( .A0(n1867), .A1(n2877), .B0(n1844), .Y(n1845) );
  AOI22XL U1841 ( .A0(n1859), .A1(x[28]), .B0(n1854), .B1(x[34]), .Y(n1832) );
  NAND2X1 U1842 ( .A(n1828), .B(n1827), .Y(n2512) );
  AOI22XL U1843 ( .A0(n2721), .A1(n1816), .B0(n1916), .B1(x[72]), .Y(n1828) );
  AOI22XL U1844 ( .A0(n2714), .A1(n1826), .B0(n2681), .B1(n1825), .Y(n1827) );
  NAND4XL U1845 ( .A(n1815), .B(n1814), .C(n1813), .D(n1812), .Y(n1816) );
  AOI211XL U1846 ( .A0(n1978), .A1(y[55]), .B0(n2003), .C0(n2002), .Y(n2230)
         );
  AOI22XL U1847 ( .A0(n2903), .A1(n1759), .B0(x[54]), .B1(n1758), .Y(n1999) );
  AOI22XL U1848 ( .A0(y[29]), .A1(n2248), .B0(y[35]), .B1(n2249), .Y(n2045) );
  AOI22XL U1849 ( .A0(y[20]), .A1(n2244), .B0(y[23]), .B1(n2245), .Y(n2047) );
  AOI22XL U1850 ( .A0(y[14]), .A1(n2242), .B0(y[17]), .B1(n2243), .Y(n2048) );
  AOI211XL U1851 ( .A0(n1978), .A1(y[58]), .B0(n1992), .C0(n1991), .Y(n1993)
         );
  INVX1 U1852 ( .A(n1910), .Y(n2515) );
  AOI211XL U1853 ( .A0(n1978), .A1(y[49]), .B0(n1998), .C0(n1997), .Y(n2237)
         );
  AOI22XL U1854 ( .A0(n2882), .A1(n1759), .B0(x[48]), .B1(n1758), .Y(n1994) );
  AOI211XL U1855 ( .A0(n1978), .A1(y[46]), .B0(n1988), .C0(n1987), .Y(n2236)
         );
  AOI22XL U1856 ( .A0(n2885), .A1(n1759), .B0(x[45]), .B1(n1758), .Y(n1984) );
  OAI2BB2XL U1857 ( .B0(y[59]), .B1(n2231), .A0N(n2907), .A1N(n2230), .Y(n2241) );
  NAND2X1 U1858 ( .A(n1791), .B(n1790), .Y(n2518) );
  AOI22XL U1859 ( .A0(n1916), .A1(y[73]), .B0(n2681), .B1(n1777), .Y(n1791) );
  AOI22XL U1860 ( .A0(n2714), .A1(n1789), .B0(n2721), .B1(n1788), .Y(n1790) );
  NAND4XL U1861 ( .A(n1776), .B(n1775), .C(n1774), .D(n1773), .Y(n1777) );
  AOI22XL U1862 ( .A0(n1916), .A1(y[74]), .B0(n2681), .B1(n1915), .Y(n1928) );
  AOI22XL U1863 ( .A0(n2714), .A1(n1926), .B0(n2721), .B1(n1925), .Y(n1927) );
  NAND4XL U1864 ( .A(n1914), .B(n1913), .C(n1912), .D(n1911), .Y(n1915) );
  NAND2X2 U1865 ( .A(n1769), .B(n2591), .Y(n2628) );
  AOI211XL U1866 ( .A0(n1978), .A1(y[31]), .B0(n2034), .C0(n2033), .Y(n2247)
         );
  AOI22XL U1867 ( .A0(n2900), .A1(n1759), .B0(x[30]), .B1(n1758), .Y(n2030) );
  AOI211XL U1868 ( .A0(n1978), .A1(y[25]), .B0(n2029), .C0(n2028), .Y(n2246)
         );
  AOI22XL U1869 ( .A0(n2889), .A1(n1759), .B0(x[24]), .B1(n1758), .Y(n2025) );
  NOR2X1 U1870 ( .A(in_valid), .B(n2670), .Y(n2675) );
  NAND4XL U1871 ( .A(n1853), .B(n1852), .C(n1851), .D(n1850), .Y(n1869) );
  OAI21XL U1872 ( .A0(n1867), .A1(n2880), .B0(n1866), .Y(n1868) );
  AOI22XL U1873 ( .A0(n1859), .A1(x[29]), .B0(n1765), .B1(x[35]), .Y(n1852) );
  AOI221XL U1874 ( .A0(x[40]), .A1(n1968), .B0(x[41]), .B1(n1757), .C0(n1969), 
        .Y(n1970) );
  OAI22XL U1875 ( .A0(x[40]), .A1(n1968), .B0(n2798), .B1(x[41]), .Y(n1969) );
  AOI221XL U1876 ( .A0(x[37]), .A1(n1968), .B0(x[38]), .B1(n1757), .C0(n1963), 
        .Y(n1964) );
  OAI22XL U1877 ( .A0(x[37]), .A1(n1968), .B0(n1757), .B1(x[38]), .Y(n1963) );
  AOI221XL U1878 ( .A0(x[43]), .A1(n1968), .B0(x[44]), .B1(n1757), .C0(n1974), 
        .Y(n1975) );
  OAI22XL U1879 ( .A0(x[43]), .A1(n1968), .B0(n2798), .B1(x[44]), .Y(n1974) );
  AOI221XL U1880 ( .A0(x[53]), .A1(n1757), .B0(n1968), .B1(x[52]), .C0(n1980), 
        .Y(n1981) );
  OAI22XL U1881 ( .A0(x[53]), .A1(n1757), .B0(x[52]), .B1(n1968), .Y(n1980) );
  AOI22XL U1882 ( .A0(y[26]), .A1(n2246), .B0(y[32]), .B1(n2247), .Y(n2046) );
  AOI221XL U1883 ( .A0(x[61]), .A1(n1968), .B0(x[62]), .B1(n1757), .C0(n1951), 
        .Y(n1952) );
  OAI22XL U1884 ( .A0(x[61]), .A1(n1968), .B0(n1757), .B1(x[62]), .Y(n1951) );
  AOI221XL U1885 ( .A0(x[64]), .A1(n1968), .B0(x[65]), .B1(n1757), .C0(n1956), 
        .Y(n1957) );
  OAI22XL U1886 ( .A0(x[64]), .A1(n1968), .B0(n1757), .B1(x[65]), .Y(n1956) );
  AOI22XL U1887 ( .A0(x[73]), .A1(n1968), .B0(n2880), .B1(n1764), .Y(n1945) );
  AOI22XL U1888 ( .A0(n2886), .A1(n1759), .B0(x[72]), .B1(n1758), .Y(n1946) );
  AOI221XL U1889 ( .A0(x[1]), .A1(n1968), .B0(x[2]), .B1(n1757), .C0(n1886), 
        .Y(n1887) );
  OAI22XL U1890 ( .A0(x[1]), .A1(n1968), .B0(n2798), .B1(x[2]), .Y(n1886) );
  AOI22XL U1891 ( .A0(x[11]), .A1(n1757), .B0(x[10]), .B1(n1968), .Y(n1895) );
  AOI22XL U1892 ( .A0(n2881), .A1(n1759), .B0(x[9]), .B1(n1758), .Y(n1896) );
  AOI22XL U1893 ( .A0(x[5]), .A1(n1757), .B0(x[4]), .B1(n1968), .Y(n1900) );
  AOI22XL U1894 ( .A0(n2894), .A1(n1759), .B0(x[3]), .B1(n1758), .Y(n1901) );
  INVX1 U1895 ( .A(n2518), .Y(n1933) );
  AOI211XL U1896 ( .A0(n1978), .A1(y[22]), .B0(n2024), .C0(n2023), .Y(n2245)
         );
  AOI22XL U1897 ( .A0(n2884), .A1(n1759), .B0(x[21]), .B1(n1758), .Y(n2020) );
  AOI211XL U1898 ( .A0(n1978), .A1(y[19]), .B0(n2019), .C0(n2018), .Y(n2244)
         );
  AOI22XL U1899 ( .A0(n2899), .A1(n1759), .B0(x[18]), .B1(n1758), .Y(n2015) );
  AOI211XL U1900 ( .A0(n1978), .A1(y[16]), .B0(n2014), .C0(n2013), .Y(n2243)
         );
  AOI22XL U1901 ( .A0(n2890), .A1(n1759), .B0(x[15]), .B1(n1758), .Y(n2010) );
  AOI211XL U1902 ( .A0(n1978), .A1(y[13]), .B0(n2009), .C0(n2008), .Y(n2242)
         );
  AOI22XL U1903 ( .A0(n2898), .A1(n1759), .B0(x[12]), .B1(n1758), .Y(n2005) );
  AOI211XL U1904 ( .A0(n1978), .A1(y[34]), .B0(n2044), .C0(n2043), .Y(n2249)
         );
  AOI22XL U1905 ( .A0(n2891), .A1(n1759), .B0(x[33]), .B1(n1758), .Y(n2040) );
  AOI211XL U1906 ( .A0(n1978), .A1(y[28]), .B0(n2039), .C0(n2038), .Y(n2248)
         );
  AOI22XL U1907 ( .A0(n2896), .A1(n1759), .B0(x[27]), .B1(n1758), .Y(n2035) );
  AOI22XL U1908 ( .A0(n2868), .A1(n2247), .B0(n2916), .B1(n2246), .Y(n2251) );
  XOR2XL U1909 ( .A(n1872), .B(n2521), .Y(n1847) );
  NOR2X2 U1910 ( .A(n2678), .B(n1778), .Y(n2714) );
  NOR2X2 U1911 ( .A(n1783), .B(n1778), .Y(n2681) );
  NOR2X2 U1912 ( .A(n2675), .B(n2801), .Y(n2719) );
  INVX1 U1913 ( .A(n2675), .Y(n2797) );
  AOI211XL U1914 ( .A0(y[69]), .A1(n2685), .B0(n2221), .C0(n2220), .Y(n2222)
         );
  OAI21XL U1915 ( .A0(n2912), .A1(n2214), .B0(n2213), .Y(n2215) );
  AOI2BB2XL U1916 ( .B0(y[2]), .B1(n2212), .A0N(n2906), .A1N(n2211), .Y(n2213)
         );
  OAI21XL U1917 ( .A0(n1978), .A1(y[7]), .B0(n1894), .Y(n2216) );
  AOI211XL U1918 ( .A0(n1978), .A1(y[7]), .B0(n1893), .C0(n1892), .Y(n1894) );
  AOI22XL U1919 ( .A0(n2872), .A1(n2257), .B0(n2922), .B1(n2256), .Y(n2258) );
  AOI211XL U1920 ( .A0(n1978), .A1(y[67]), .B0(n1944), .C0(n1943), .Y(n2261)
         );
  AOI22XL U1921 ( .A0(n2895), .A1(n1759), .B0(x[66]), .B1(n1758), .Y(n1940) );
  AOI22XL U1922 ( .A0(n2871), .A1(n2233), .B0(n2920), .B1(n2232), .Y(n2240) );
  AOI22XL U1923 ( .A0(n2865), .A1(n2237), .B0(n2914), .B1(n2236), .Y(n2238) );
  AOI22XL U1924 ( .A0(n2867), .A1(n2235), .B0(n2921), .B1(n2234), .Y(n2239) );
  AOI22XL U1925 ( .A0(n2870), .A1(n2249), .B0(n2917), .B1(n2248), .Y(n2250) );
  AOI22XL U1926 ( .A0(n2869), .A1(n2243), .B0(n2918), .B1(n2242), .Y(n2253) );
  AOI22XL U1927 ( .A0(n2866), .A1(n2245), .B0(n2919), .B1(n2244), .Y(n2252) );
  NAND2X1 U1928 ( .A(n2721), .B(n2720), .Y(n2789) );
  NAND2X1 U1929 ( .A(n2714), .B(n2720), .Y(n2771) );
  NAND2X1 U1930 ( .A(n2681), .B(n2720), .Y(n2758) );
  CLKINVX2 U1931 ( .A(n2719), .Y(n2760) );
  NOR2X2 U1932 ( .A(n2861), .B(n2862), .Y(n2674) );
  NAND2XL U1933 ( .A(n2853), .B(n2591), .Y(n2670) );
  OAI21XL U1934 ( .A0(n1929), .A1(n1910), .B0(n1909), .Y(n1939) );
  OAI21XL U1935 ( .A0(n1937), .A1(n2530), .B0(n1936), .Y(n1938) );
  NAND2X1 U1936 ( .A(n1766), .B(n2399), .Y(n2635) );
  NAND2XL U1937 ( .A(cnt[1]), .B(N2025), .Y(n2844) );
  INVXL U1938 ( .A(n2838), .Y(n2847) );
  NOR2X2 U1939 ( .A(in_valid), .B(n2628), .Y(n2720) );
  INVX1 U1940 ( .A(n2720), .Y(n2846) );
  NAND2XL U1941 ( .A(n2671), .B(n2670), .Y(n2838) );
  NAND2X1 U1942 ( .A(n2266), .B(n2265), .Y(n2267) );
  AOI22X1 U1943 ( .A0(n2057), .A1(n2688), .B0(n2056), .B1(n2055), .Y(n2268) );
  NOR4X1 U1944 ( .A(n2229), .B(n2274), .C(n2228), .D(n2227), .Y(n2266) );
  NOR2BXL U1945 ( .AN(n2390), .B(n2853), .Y(n2854) );
  AOI22XL U1946 ( .A0(n2738), .A1(x[13]), .B0(n1763), .B1(x[19]), .Y(n1839) );
  AOI22XL U1947 ( .A0(n1761), .A1(x[1]), .B0(n1760), .B1(x[7]), .Y(n1841) );
  AOI22XL U1948 ( .A0(n1766), .A1(x[22]), .B0(n1762), .B1(x[16]), .Y(n1838) );
  AOI22XL U1949 ( .A0(n1859), .A1(x[4]), .B0(n1854), .B1(x[10]), .Y(n1840) );
  AOI22XL U1950 ( .A0(n1761), .A1(x[49]), .B0(n1760), .B1(x[55]), .Y(n1837) );
  AOI22XL U1951 ( .A0(n1766), .A1(x[70]), .B0(n1762), .B1(x[64]), .Y(n1834) );
  AOI22XL U1952 ( .A0(n1767), .A1(x[61]), .B0(n1763), .B1(x[67]), .Y(n1835) );
  AOI22XL U1953 ( .A0(n2738), .A1(x[14]), .B0(n1763), .B1(x[20]), .Y(n1861) );
  AOI22XL U1954 ( .A0(n1761), .A1(x[2]), .B0(n1760), .B1(x[8]), .Y(n1863) );
  AOI22XL U1955 ( .A0(n1766), .A1(x[23]), .B0(n1762), .B1(x[17]), .Y(n1860) );
  AOI22XL U1956 ( .A0(n1859), .A1(x[5]), .B0(n1765), .B1(x[11]), .Y(n1862) );
  AOI22XL U1957 ( .A0(n2738), .A1(x[62]), .B0(n1763), .B1(x[68]), .Y(n1856) );
  AOI22XL U1958 ( .A0(n1761), .A1(x[50]), .B0(n1760), .B1(x[56]), .Y(n1858) );
  AOI22XL U1959 ( .A0(n1766), .A1(x[71]), .B0(n1762), .B1(x[65]), .Y(n1855) );
  AOI22XL U1960 ( .A0(n1761), .A1(x[0]), .B0(n1760), .B1(x[6]), .Y(n1824) );
  AOI22XL U1961 ( .A0(n1761), .A1(x[24]), .B0(n1760), .B1(x[30]), .Y(n1820) );
  NOR2XL U1962 ( .A(direction[1]), .B(n1872), .Y(n1875) );
  NAND2XL U1963 ( .A(n1873), .B(n1878), .Y(n1874) );
  AOI2BB1XL U1964 ( .A0N(n1873), .A1N(n1878), .B0(n2512), .Y(n1870) );
  AOI22XL U1965 ( .A0(direction[2]), .A1(n2521), .B0(n1878), .B1(n2878), .Y(
        n1880) );
  AOI221XL U1966 ( .A0(x[31]), .A1(n1968), .B0(x[32]), .B1(n1757), .C0(n2031), 
        .Y(n2032) );
  OAI22XL U1967 ( .A0(x[31]), .A1(n1968), .B0(n2798), .B1(x[32]), .Y(n2031) );
  AOI221XL U1968 ( .A0(x[25]), .A1(n1968), .B0(x[26]), .B1(n1757), .C0(n2026), 
        .Y(n2027) );
  OAI22XL U1969 ( .A0(x[25]), .A1(n1968), .B0(n2798), .B1(x[26]), .Y(n2026) );
  AOI22XL U1970 ( .A0(n2496), .A1(n2447), .B0(n2509), .B1(n2446), .Y(n2448) );
  NAND4XL U1971 ( .A(n2441), .B(n2440), .C(n2439), .D(n2438), .Y(n2447) );
  NAND4XL U1972 ( .A(n2445), .B(n2444), .C(n2443), .D(n2442), .Y(n2446) );
  AOI22XL U1973 ( .A0(n2721), .A1(n1843), .B0(n2681), .B1(n1842), .Y(n1844) );
  NAND4XL U1974 ( .A(n1837), .B(n1836), .C(n1835), .D(n1834), .Y(n1843) );
  NAND4XL U1975 ( .A(n1841), .B(n1840), .C(n1839), .D(n1838), .Y(n1842) );
  AOI22XL U1976 ( .A0(n1859), .A1(x[52]), .B0(n1854), .B1(x[58]), .Y(n1836) );
  AOI22XL U1977 ( .A0(n1761), .A1(x[25]), .B0(n1760), .B1(x[31]), .Y(n1833) );
  AOI22XL U1978 ( .A0(n1766), .A1(x[46]), .B0(n1762), .B1(x[40]), .Y(n1830) );
  AOI22XL U1979 ( .A0(n1767), .A1(x[37]), .B0(n1763), .B1(x[43]), .Y(n1831) );
  AOI22XL U1980 ( .A0(n2721), .A1(n1865), .B0(n2681), .B1(n1864), .Y(n1866) );
  NAND4XL U1981 ( .A(n1858), .B(n1857), .C(n1856), .D(n1855), .Y(n1865) );
  NAND4XL U1982 ( .A(n1863), .B(n1862), .C(n1861), .D(n1860), .Y(n1864) );
  AOI22XL U1983 ( .A0(n1859), .A1(x[53]), .B0(n1854), .B1(x[59]), .Y(n1857) );
  AOI22XL U1984 ( .A0(n2738), .A1(x[38]), .B0(n1763), .B1(x[44]), .Y(n1851) );
  AOI22XL U1985 ( .A0(n1761), .A1(x[26]), .B0(n1760), .B1(x[32]), .Y(n1853) );
  AOI22XL U1986 ( .A0(n1766), .A1(x[47]), .B0(n1762), .B1(x[41]), .Y(n1850) );
  AOI22XL U1987 ( .A0(n2394), .A1(n2861), .B0(cnt[3]), .B1(n2393), .Y(n2407)
         );
  AOI22XL U1988 ( .A0(n1761), .A1(x[48]), .B0(n1760), .B1(x[54]), .Y(n1815) );
  AOI22XL U1989 ( .A0(n1766), .A1(x[69]), .B0(n1762), .B1(x[63]), .Y(n1812) );
  AOI22XL U1990 ( .A0(n1767), .A1(x[60]), .B0(n1763), .B1(x[66]), .Y(n1813) );
  AOI22XL U1991 ( .A0(n1859), .A1(x[51]), .B0(n1854), .B1(x[57]), .Y(n1814) );
  NAND4XL U1992 ( .A(n1824), .B(n1823), .C(n1822), .D(n1821), .Y(n1825) );
  AOI22XL U1993 ( .A0(n1859), .A1(x[3]), .B0(n1854), .B1(x[9]), .Y(n1823) );
  AOI22XL U1994 ( .A0(n1767), .A1(x[12]), .B0(n1763), .B1(x[18]), .Y(n1822) );
  AOI22XL U1995 ( .A0(n1766), .A1(x[21]), .B0(n1762), .B1(x[15]), .Y(n1821) );
  NAND4XL U1996 ( .A(n1820), .B(n1819), .C(n1818), .D(n1817), .Y(n1826) );
  AOI22XL U1997 ( .A0(n1859), .A1(x[27]), .B0(n1854), .B1(x[33]), .Y(n1819) );
  AOI22XL U1998 ( .A0(n1767), .A1(x[36]), .B0(n1763), .B1(x[42]), .Y(n1818) );
  AOI22XL U1999 ( .A0(n1766), .A1(x[45]), .B0(n1762), .B1(x[39]), .Y(n1817) );
  AOI22XL U2000 ( .A0(n2496), .A1(n2486), .B0(n2507), .B1(n2485), .Y(n2487) );
  NAND4XL U2001 ( .A(n2480), .B(n2479), .C(n2478), .D(n2477), .Y(n2486) );
  NAND4XL U2002 ( .A(n2484), .B(n2483), .C(n2482), .D(n2481), .Y(n2485) );
  NAND4XL U2003 ( .A(n2420), .B(n2419), .C(n2418), .D(n2417), .Y(n2421) );
  NAND4XL U2004 ( .A(n2429), .B(n2428), .C(n2427), .D(n2426), .Y(n2430) );
  INVXL U2005 ( .A(n2407), .Y(n2400) );
  NAND2BXL U2006 ( .AN(n2399), .B(n2401), .Y(n2406) );
  AOI22XL U2007 ( .A0(n2743), .A1(have_tried_direction[128]), .B0(n2750), .B1(
        have_tried_direction[8]), .Y(n2197) );
  AOI22XL U2008 ( .A0(n2840), .A1(have_tried_direction[120]), .B0(n2192), .B1(
        have_tried_direction[136]), .Y(n2196) );
  AOI22XL U2009 ( .A0(n2761), .A1(have_tried_direction[16]), .B0(n2191), .B1(
        have_tried_direction[184]), .Y(n2198) );
  AOI22XL U2010 ( .A0(n2194), .A1(have_tried_direction[144]), .B0(n2193), .B1(
        have_tried_direction[152]), .Y(n2195) );
  AOI22XL U2011 ( .A0(n2703), .A1(have_tried_direction[32]), .B0(n2695), .B1(
        have_tried_direction[40]), .Y(n2189) );
  AOI22XL U2012 ( .A0(n2743), .A1(have_tried_direction[129]), .B0(n2750), .B1(
        have_tried_direction[9]), .Y(n2168) );
  AOI22XL U2013 ( .A0(n2840), .A1(have_tried_direction[121]), .B0(n2192), .B1(
        have_tried_direction[137]), .Y(n2167) );
  AOI22XL U2014 ( .A0(n2761), .A1(have_tried_direction[17]), .B0(n2191), .B1(
        have_tried_direction[185]), .Y(n2169) );
  AOI22XL U2015 ( .A0(n2194), .A1(have_tried_direction[145]), .B0(n2193), .B1(
        have_tried_direction[153]), .Y(n2166) );
  AOI22XL U2016 ( .A0(n2703), .A1(have_tried_direction[33]), .B0(n2695), .B1(
        have_tried_direction[41]), .Y(n2164) );
  AOI22XL U2017 ( .A0(n2743), .A1(have_tried_direction[130]), .B0(n2750), .B1(
        have_tried_direction[10]), .Y(n2152) );
  AOI22XL U2018 ( .A0(n2840), .A1(have_tried_direction[122]), .B0(n2192), .B1(
        have_tried_direction[138]), .Y(n2151) );
  AOI22XL U2019 ( .A0(n2761), .A1(have_tried_direction[18]), .B0(n2191), .B1(
        have_tried_direction[186]), .Y(n2153) );
  AOI22XL U2020 ( .A0(n2194), .A1(have_tried_direction[146]), .B0(n2193), .B1(
        have_tried_direction[154]), .Y(n2150) );
  AOI22XL U2021 ( .A0(n2703), .A1(have_tried_direction[34]), .B0(n2695), .B1(
        have_tried_direction[42]), .Y(n2148) );
  AOI22XL U2022 ( .A0(n2743), .A1(have_tried_direction[131]), .B0(n2750), .B1(
        have_tried_direction[11]), .Y(n2136) );
  AOI22XL U2023 ( .A0(n2840), .A1(have_tried_direction[123]), .B0(n2192), .B1(
        have_tried_direction[139]), .Y(n2135) );
  AOI22XL U2024 ( .A0(n2761), .A1(have_tried_direction[19]), .B0(n2191), .B1(
        have_tried_direction[187]), .Y(n2137) );
  AOI22XL U2025 ( .A0(n2194), .A1(have_tried_direction[147]), .B0(n2193), .B1(
        have_tried_direction[155]), .Y(n2134) );
  AOI22XL U2026 ( .A0(n2703), .A1(have_tried_direction[35]), .B0(n2695), .B1(
        have_tried_direction[43]), .Y(n2132) );
  AOI22XL U2027 ( .A0(n2743), .A1(have_tried_direction[132]), .B0(n2750), .B1(
        have_tried_direction[12]), .Y(n2116) );
  AOI22XL U2028 ( .A0(n2840), .A1(have_tried_direction[124]), .B0(n2192), .B1(
        have_tried_direction[140]), .Y(n2115) );
  AOI22XL U2029 ( .A0(n2761), .A1(have_tried_direction[20]), .B0(n2191), .B1(
        have_tried_direction[188]), .Y(n2117) );
  AOI22XL U2030 ( .A0(n2194), .A1(have_tried_direction[148]), .B0(n2193), .B1(
        have_tried_direction[156]), .Y(n2114) );
  AOI22XL U2031 ( .A0(n2703), .A1(have_tried_direction[36]), .B0(n2695), .B1(
        have_tried_direction[44]), .Y(n2112) );
  AOI22XL U2032 ( .A0(n2743), .A1(have_tried_direction[133]), .B0(n2750), .B1(
        have_tried_direction[13]), .Y(n2100) );
  AOI22XL U2033 ( .A0(n2840), .A1(have_tried_direction[125]), .B0(n2192), .B1(
        have_tried_direction[141]), .Y(n2099) );
  AOI22XL U2034 ( .A0(n2761), .A1(have_tried_direction[21]), .B0(n2191), .B1(
        have_tried_direction[189]), .Y(n2101) );
  AOI22XL U2035 ( .A0(n2194), .A1(have_tried_direction[149]), .B0(n2193), .B1(
        have_tried_direction[157]), .Y(n2098) );
  AOI22XL U2036 ( .A0(n2703), .A1(have_tried_direction[37]), .B0(n2695), .B1(
        have_tried_direction[45]), .Y(n2096) );
  AOI22XL U2037 ( .A0(n2743), .A1(have_tried_direction[134]), .B0(n2750), .B1(
        have_tried_direction[14]), .Y(n2084) );
  AOI22XL U2038 ( .A0(n2840), .A1(have_tried_direction[126]), .B0(n2192), .B1(
        have_tried_direction[142]), .Y(n2083) );
  AOI22XL U2039 ( .A0(n2761), .A1(have_tried_direction[22]), .B0(n2191), .B1(
        have_tried_direction[190]), .Y(n2085) );
  AOI22XL U2040 ( .A0(n2194), .A1(have_tried_direction[150]), .B0(n2193), .B1(
        have_tried_direction[158]), .Y(n2082) );
  AOI22XL U2041 ( .A0(n2703), .A1(have_tried_direction[38]), .B0(n2695), .B1(
        have_tried_direction[46]), .Y(n2080) );
  AOI221XL U2042 ( .A0(x[55]), .A1(n1968), .B0(x[56]), .B1(n1757), .C0(n2000), 
        .Y(n2001) );
  OAI22XL U2043 ( .A0(x[55]), .A1(n1968), .B0(n2798), .B1(x[56]), .Y(n2000) );
  AOI22XL U2044 ( .A0(x[59]), .A1(n1757), .B0(x[58]), .B1(n1968), .Y(n1989) );
  AOI22XL U2045 ( .A0(n2893), .A1(n1759), .B0(x[57]), .B1(n1758), .Y(n1990) );
  AOI22XL U2046 ( .A0(n2738), .A1(y[37]), .B0(n1763), .B1(y[43]), .Y(n1780) );
  AOI22XL U2047 ( .A0(n1761), .A1(y[49]), .B0(n1760), .B1(y[55]), .Y(n1787) );
  AOI22XL U2048 ( .A0(n2738), .A1(y[62]), .B0(n1763), .B1(y[68]), .Y(n1922) );
  AOI22XL U2049 ( .A0(n2738), .A1(y[38]), .B0(n1763), .B1(y[44]), .Y(n1918) );
  AOI22XL U2050 ( .A0(n1761), .A1(y[48]), .B0(n1760), .B1(y[54]), .Y(n1804) );
  AOI22XL U2051 ( .A0(n1766), .A1(y[45]), .B0(n1762), .B1(y[39]), .Y(n1797) );
  AOI221XL U2052 ( .A0(x[49]), .A1(n1968), .B0(x[50]), .B1(n1757), .C0(n1995), 
        .Y(n1996) );
  OAI22XL U2053 ( .A0(x[49]), .A1(n1968), .B0(n2798), .B1(x[50]), .Y(n1995) );
  AOI221XL U2054 ( .A0(x[46]), .A1(n1968), .B0(x[47]), .B1(n1757), .C0(n1985), 
        .Y(n1986) );
  OAI22XL U2055 ( .A0(x[46]), .A1(n1968), .B0(n2798), .B1(x[47]), .Y(n1985) );
  AOI221XL U2056 ( .A0(x[22]), .A1(n1968), .B0(x[23]), .B1(n1757), .C0(n2021), 
        .Y(n2022) );
  OAI22XL U2057 ( .A0(x[22]), .A1(n1968), .B0(n2798), .B1(x[23]), .Y(n2021) );
  AOI221XL U2058 ( .A0(x[19]), .A1(n1968), .B0(x[20]), .B1(n1757), .C0(n2016), 
        .Y(n2017) );
  OAI22XL U2059 ( .A0(x[19]), .A1(n1968), .B0(n2798), .B1(x[20]), .Y(n2016) );
  AOI221XL U2060 ( .A0(x[16]), .A1(n1968), .B0(x[17]), .B1(n1757), .C0(n2011), 
        .Y(n2012) );
  OAI22XL U2061 ( .A0(x[16]), .A1(n1968), .B0(n2798), .B1(x[17]), .Y(n2011) );
  AOI221XL U2062 ( .A0(x[13]), .A1(n1968), .B0(x[14]), .B1(n1757), .C0(n2006), 
        .Y(n2007) );
  OAI22XL U2063 ( .A0(x[13]), .A1(n1968), .B0(n2798), .B1(x[14]), .Y(n2006) );
  AOI221XL U2064 ( .A0(x[34]), .A1(n1968), .B0(x[35]), .B1(n1757), .C0(n2041), 
        .Y(n2042) );
  OAI22XL U2065 ( .A0(x[34]), .A1(n1968), .B0(n2798), .B1(x[35]), .Y(n2041) );
  AOI221XL U2066 ( .A0(x[28]), .A1(n1968), .B0(x[29]), .B1(n1757), .C0(n2036), 
        .Y(n2037) );
  OAI22XL U2067 ( .A0(x[28]), .A1(n1968), .B0(n1757), .B1(x[29]), .Y(n2036) );
  NOR2XL U2068 ( .A(n2592), .B(n2588), .Y(n1877) );
  INVX1 U2069 ( .A(n2678), .Y(n1783) );
  NAND4XL U2070 ( .A(n2437), .B(n2436), .C(n2435), .D(n2434), .Y(n2450) );
  NAND4XL U2071 ( .A(n2494), .B(n2493), .C(n2492), .D(n2491), .Y(n2495) );
  NAND4XL U2072 ( .A(n2505), .B(n2504), .C(n2503), .D(n2502), .Y(n2506) );
  NAND4XL U2073 ( .A(n2501), .B(n2500), .C(n2499), .D(n2498), .Y(n2508) );
  NOR2X1 U2074 ( .A(n2407), .B(n2406), .Y(n2509) );
  NAND4XL U2075 ( .A(n2468), .B(n2467), .C(n2466), .D(n2465), .Y(n2469) );
  NAND4XL U2076 ( .A(n2464), .B(n2463), .C(n2462), .D(n2461), .Y(n2470) );
  NAND4XL U2077 ( .A(n2459), .B(n2458), .C(n2457), .D(n2456), .Y(n2460) );
  INVXL U2078 ( .A(n2488), .Y(n2497) );
  AOI21XL U2079 ( .A0(n2509), .A1(n2490), .B0(n2489), .Y(n2513) );
  NAND4XL U2080 ( .A(n2476), .B(n2475), .C(n2474), .D(n2473), .Y(n2490) );
  NOR2XL U2081 ( .A(n2513), .B(n2512), .Y(n2520) );
  NAND2XL U2082 ( .A(n2433), .B(n2432), .Y(n2514) );
  AOI22XL U2083 ( .A0(n2509), .A1(n2431), .B0(n2496), .B1(n2430), .Y(n2432) );
  AOI22XL U2084 ( .A0(y[72]), .A1(n2497), .B0(n2507), .B1(n2421), .Y(n2433) );
  NAND4XL U2085 ( .A(n2425), .B(n2424), .C(n2423), .D(n2422), .Y(n2431) );
  AOI22XL U2086 ( .A0(n2496), .A1(n2413), .B0(n2509), .B1(n2412), .Y(n2414) );
  NAND4XL U2087 ( .A(n2405), .B(n2404), .C(n2403), .D(n2402), .Y(n2413) );
  NAND4XL U2088 ( .A(n2411), .B(n2410), .C(n2409), .D(n2408), .Y(n2412) );
  NAND2XL U2089 ( .A(n2406), .B(n2400), .Y(n2488) );
  NAND2XL U2090 ( .A(n2515), .B(n2514), .Y(n2516) );
  AOI22XL U2091 ( .A0(x[71]), .A1(n1757), .B0(y[70]), .B1(n1978), .Y(n2217) );
  AOI22XL U2092 ( .A0(x[70]), .A1(n1968), .B0(n2219), .B1(n2905), .Y(n2218) );
  AOI21XL U2093 ( .A0(n1933), .A1(n2879), .B0(n1810), .Y(n1811) );
  XOR2XL U2094 ( .A(n1933), .B(n2515), .Y(n1809) );
  AOI22XL U2095 ( .A0(n2743), .A1(have_tried_direction[135]), .B0(n2750), .B1(
        have_tried_direction[15]), .Y(n2068) );
  AOI22XL U2096 ( .A0(n2840), .A1(have_tried_direction[127]), .B0(n2192), .B1(
        have_tried_direction[143]), .Y(n2067) );
  AOI22XL U2097 ( .A0(n2761), .A1(have_tried_direction[23]), .B0(n2191), .B1(
        have_tried_direction[191]), .Y(n2069) );
  AOI22XL U2098 ( .A0(n2194), .A1(have_tried_direction[151]), .B0(n2193), .B1(
        have_tried_direction[159]), .Y(n2066) );
  AOI22XL U2099 ( .A0(n2703), .A1(have_tried_direction[39]), .B0(n2695), .B1(
        have_tried_direction[47]), .Y(n2064) );
  AOI22XL U2100 ( .A0(n2711), .A1(have_tried_direction[63]), .B0(n2179), .B1(
        have_tried_direction[87]), .Y(n2062) );
  AOI22XL U2101 ( .A0(n2711), .A1(have_tried_direction[56]), .B0(n2179), .B1(
        have_tried_direction[80]), .Y(n2188) );
  AOI22XL U2102 ( .A0(n2183), .A1(have_tried_direction[72]), .B0(n2182), .B1(
        have_tried_direction[96]), .Y(n2186) );
  AOI22XL U2103 ( .A0(n2699), .A1(have_tried_direction[0]), .B0(n2184), .B1(
        have_tried_direction[104]), .Y(n2185) );
  AOI22XL U2104 ( .A0(n2181), .A1(have_tried_direction[88]), .B0(n2180), .B1(
        have_tried_direction[112]), .Y(n2187) );
  AOI211XL U2105 ( .A0(n2707), .A1(have_tried_direction[48]), .B0(n2200), .C0(
        n2199), .Y(n2201) );
  NAND2XL U2106 ( .A(n2190), .B(n2189), .Y(n2200) );
  NAND4XL U2107 ( .A(n2198), .B(n2197), .C(n2196), .D(n2195), .Y(n2199) );
  AOI22XL U2108 ( .A0(n2674), .A1(have_tried_direction[192]), .B0(n2755), .B1(
        have_tried_direction[64]), .Y(n2190) );
  AOI22XL U2109 ( .A0(n2711), .A1(have_tried_direction[57]), .B0(n2179), .B1(
        have_tried_direction[81]), .Y(n2163) );
  AOI22XL U2110 ( .A0(n2183), .A1(have_tried_direction[73]), .B0(n2182), .B1(
        have_tried_direction[97]), .Y(n2161) );
  AOI22XL U2111 ( .A0(n2699), .A1(have_tried_direction[1]), .B0(n2184), .B1(
        have_tried_direction[105]), .Y(n2160) );
  AOI22XL U2112 ( .A0(n2181), .A1(have_tried_direction[89]), .B0(n2180), .B1(
        have_tried_direction[113]), .Y(n2162) );
  AOI211XL U2113 ( .A0(n2707), .A1(have_tried_direction[49]), .B0(n2171), .C0(
        n2170), .Y(n2172) );
  NAND2XL U2114 ( .A(n2165), .B(n2164), .Y(n2171) );
  NAND4XL U2115 ( .A(n2169), .B(n2168), .C(n2167), .D(n2166), .Y(n2170) );
  AOI22XL U2116 ( .A0(n2674), .A1(have_tried_direction[193]), .B0(n2755), .B1(
        have_tried_direction[65]), .Y(n2165) );
  AOI22XL U2117 ( .A0(n2711), .A1(have_tried_direction[58]), .B0(n2179), .B1(
        have_tried_direction[82]), .Y(n2147) );
  AOI22XL U2118 ( .A0(n2183), .A1(have_tried_direction[74]), .B0(n2182), .B1(
        have_tried_direction[98]), .Y(n2145) );
  AOI22XL U2119 ( .A0(n2699), .A1(have_tried_direction[2]), .B0(n2184), .B1(
        have_tried_direction[106]), .Y(n2144) );
  AOI22XL U2120 ( .A0(n2181), .A1(have_tried_direction[90]), .B0(n2180), .B1(
        have_tried_direction[114]), .Y(n2146) );
  AOI211XL U2121 ( .A0(n2707), .A1(have_tried_direction[50]), .B0(n2155), .C0(
        n2154), .Y(n2156) );
  NAND2XL U2122 ( .A(n2149), .B(n2148), .Y(n2155) );
  NAND4XL U2123 ( .A(n2153), .B(n2152), .C(n2151), .D(n2150), .Y(n2154) );
  AOI22XL U2124 ( .A0(n2674), .A1(have_tried_direction[194]), .B0(n2755), .B1(
        have_tried_direction[66]), .Y(n2149) );
  AOI22XL U2125 ( .A0(n2711), .A1(have_tried_direction[59]), .B0(n2179), .B1(
        have_tried_direction[83]), .Y(n2131) );
  AOI22XL U2126 ( .A0(n2183), .A1(have_tried_direction[75]), .B0(n2182), .B1(
        have_tried_direction[99]), .Y(n2129) );
  AOI22XL U2127 ( .A0(n2699), .A1(have_tried_direction[3]), .B0(n2184), .B1(
        have_tried_direction[107]), .Y(n2128) );
  AOI22XL U2128 ( .A0(n2181), .A1(have_tried_direction[91]), .B0(n2180), .B1(
        have_tried_direction[115]), .Y(n2130) );
  AOI211XL U2129 ( .A0(n2707), .A1(have_tried_direction[51]), .B0(n2139), .C0(
        n2138), .Y(n2140) );
  NAND2XL U2130 ( .A(n2133), .B(n2132), .Y(n2139) );
  NAND4XL U2131 ( .A(n2137), .B(n2136), .C(n2135), .D(n2134), .Y(n2138) );
  AOI22XL U2132 ( .A0(n2674), .A1(have_tried_direction[195]), .B0(n2755), .B1(
        have_tried_direction[67]), .Y(n2133) );
  AOI22XL U2133 ( .A0(n2711), .A1(have_tried_direction[60]), .B0(n2179), .B1(
        have_tried_direction[84]), .Y(n2111) );
  AOI22XL U2134 ( .A0(n2183), .A1(have_tried_direction[76]), .B0(n2182), .B1(
        have_tried_direction[100]), .Y(n2109) );
  AOI22XL U2135 ( .A0(n2699), .A1(have_tried_direction[4]), .B0(n2184), .B1(
        have_tried_direction[108]), .Y(n2108) );
  AOI22XL U2136 ( .A0(n2181), .A1(have_tried_direction[92]), .B0(n2180), .B1(
        have_tried_direction[116]), .Y(n2110) );
  AOI211XL U2137 ( .A0(n2707), .A1(have_tried_direction[52]), .B0(n2119), .C0(
        n2118), .Y(n2120) );
  NAND2XL U2138 ( .A(n2113), .B(n2112), .Y(n2119) );
  NAND4XL U2139 ( .A(n2117), .B(n2116), .C(n2115), .D(n2114), .Y(n2118) );
  AOI22XL U2140 ( .A0(n2674), .A1(have_tried_direction[196]), .B0(n2755), .B1(
        have_tried_direction[68]), .Y(n2113) );
  AOI22XL U2141 ( .A0(n2711), .A1(have_tried_direction[61]), .B0(n2179), .B1(
        have_tried_direction[85]), .Y(n2095) );
  AOI22XL U2142 ( .A0(n2183), .A1(have_tried_direction[77]), .B0(n2182), .B1(
        have_tried_direction[101]), .Y(n2093) );
  AOI22XL U2143 ( .A0(n2699), .A1(have_tried_direction[5]), .B0(n2184), .B1(
        have_tried_direction[109]), .Y(n2092) );
  AOI22XL U2144 ( .A0(n2181), .A1(have_tried_direction[93]), .B0(n2180), .B1(
        have_tried_direction[117]), .Y(n2094) );
  AOI211XL U2145 ( .A0(n2707), .A1(have_tried_direction[53]), .B0(n2103), .C0(
        n2102), .Y(n2104) );
  NAND2XL U2146 ( .A(n2097), .B(n2096), .Y(n2103) );
  NAND4XL U2147 ( .A(n2101), .B(n2100), .C(n2099), .D(n2098), .Y(n2102) );
  AOI22XL U2148 ( .A0(n2674), .A1(have_tried_direction[197]), .B0(n2755), .B1(
        have_tried_direction[69]), .Y(n2097) );
  AOI22XL U2149 ( .A0(n2711), .A1(have_tried_direction[62]), .B0(n2179), .B1(
        have_tried_direction[86]), .Y(n2079) );
  AOI22XL U2150 ( .A0(n2183), .A1(have_tried_direction[78]), .B0(n2182), .B1(
        have_tried_direction[102]), .Y(n2077) );
  AOI22XL U2151 ( .A0(n2699), .A1(have_tried_direction[6]), .B0(n2184), .B1(
        have_tried_direction[110]), .Y(n2076) );
  AOI22XL U2152 ( .A0(n2181), .A1(have_tried_direction[94]), .B0(n2180), .B1(
        have_tried_direction[118]), .Y(n2078) );
  INVX1 U2153 ( .A(n2178), .Y(n1768) );
  AOI211XL U2154 ( .A0(n2707), .A1(have_tried_direction[54]), .B0(n2087), .C0(
        n2086), .Y(n2088) );
  NAND2XL U2155 ( .A(n2081), .B(n2080), .Y(n2087) );
  NAND4XL U2156 ( .A(n2085), .B(n2084), .C(n2083), .D(n2082), .Y(n2086) );
  AOI22XL U2157 ( .A0(n2674), .A1(have_tried_direction[198]), .B0(n2755), .B1(
        have_tried_direction[70]), .Y(n2081) );
  AOI22XL U2158 ( .A0(x[8]), .A1(n1757), .B0(x[7]), .B1(n1968), .Y(n1890) );
  AOI22XL U2159 ( .A0(n2897), .A1(n1759), .B0(x[6]), .B1(n1758), .Y(n1891) );
  AOI22XL U2160 ( .A0(n2738), .A1(y[13]), .B0(n1763), .B1(y[19]), .Y(n1774) );
  AOI22XL U2161 ( .A0(n1761), .A1(y[1]), .B0(n1760), .B1(y[7]), .Y(n1776) );
  AOI22XL U2162 ( .A0(n1766), .A1(y[22]), .B0(n1762), .B1(y[16]), .Y(n1773) );
  AOI22XL U2163 ( .A0(n2765), .A1(y[4]), .B0(n1854), .B1(y[10]), .Y(n1775) );
  NAND4XL U2164 ( .A(n1782), .B(n1781), .C(n1780), .D(n1779), .Y(n1789) );
  AOI22XL U2165 ( .A0(n2765), .A1(y[28]), .B0(n1854), .B1(y[34]), .Y(n1781) );
  AOI22XL U2166 ( .A0(n1761), .A1(y[25]), .B0(n2058), .B1(y[31]), .Y(n1782) );
  AOI22XL U2167 ( .A0(n1766), .A1(y[46]), .B0(n1762), .B1(y[40]), .Y(n1779) );
  NAND4XL U2168 ( .A(n1787), .B(n1786), .C(n1785), .D(n1784), .Y(n1788) );
  AOI22XL U2169 ( .A0(n1859), .A1(y[52]), .B0(n1854), .B1(y[58]), .Y(n1786) );
  AOI22XL U2170 ( .A0(n1767), .A1(y[61]), .B0(n1763), .B1(y[67]), .Y(n1785) );
  AOI22XL U2171 ( .A0(n1766), .A1(y[70]), .B0(n1762), .B1(y[64]), .Y(n1784) );
  AOI22XL U2172 ( .A0(n2738), .A1(y[14]), .B0(n1763), .B1(y[20]), .Y(n1912) );
  AOI22XL U2173 ( .A0(n1761), .A1(y[2]), .B0(n1760), .B1(y[8]), .Y(n1914) );
  AOI22XL U2174 ( .A0(n1766), .A1(y[23]), .B0(n1762), .B1(y[17]), .Y(n1911) );
  AOI22XL U2175 ( .A0(n2765), .A1(y[5]), .B0(n1765), .B1(y[11]), .Y(n1913) );
  NAND4XL U2176 ( .A(n1924), .B(n1923), .C(n1922), .D(n1921), .Y(n1925) );
  AOI22XL U2177 ( .A0(n2765), .A1(y[53]), .B0(n1765), .B1(y[59]), .Y(n1923) );
  AOI22XL U2178 ( .A0(n1766), .A1(y[71]), .B0(n1762), .B1(y[65]), .Y(n1921) );
  AOI22XL U2179 ( .A0(n1761), .A1(y[50]), .B0(n1760), .B1(y[56]), .Y(n1924) );
  NAND4XL U2180 ( .A(n1920), .B(n1919), .C(n1918), .D(n1917), .Y(n1926) );
  AOI22XL U2181 ( .A0(n2765), .A1(y[29]), .B0(n1765), .B1(y[35]), .Y(n1919) );
  AOI22XL U2182 ( .A0(n1766), .A1(y[47]), .B0(n1762), .B1(y[41]), .Y(n1917) );
  AOI22XL U2183 ( .A0(n1761), .A1(y[26]), .B0(n1760), .B1(y[32]), .Y(n1920) );
  AOI22XL U2184 ( .A0(n1761), .A1(y[0]), .B0(n1760), .B1(y[6]), .Y(n1795) );
  AOI22XL U2185 ( .A0(n1766), .A1(y[21]), .B0(n1762), .B1(y[15]), .Y(n1792) );
  AOI22XL U2186 ( .A0(n1767), .A1(y[12]), .B0(n1763), .B1(y[18]), .Y(n1793) );
  AOI22XL U2187 ( .A0(n1859), .A1(y[3]), .B0(n1854), .B1(y[9]), .Y(n1794) );
  NAND4XL U2188 ( .A(n1804), .B(n1803), .C(n1802), .D(n1801), .Y(n1805) );
  AOI22XL U2189 ( .A0(n1859), .A1(y[51]), .B0(n1854), .B1(y[57]), .Y(n1803) );
  AOI22XL U2190 ( .A0(n1767), .A1(y[60]), .B0(n1763), .B1(y[66]), .Y(n1802) );
  AOI22XL U2191 ( .A0(n1766), .A1(y[69]), .B0(n1762), .B1(y[63]), .Y(n1801) );
  NAND4XL U2192 ( .A(n1800), .B(n1799), .C(n1798), .D(n1797), .Y(n1806) );
  AOI22XL U2193 ( .A0(n1859), .A1(y[27]), .B0(n1854), .B1(y[33]), .Y(n1799) );
  AOI22XL U2194 ( .A0(n1767), .A1(y[36]), .B0(n1763), .B1(y[42]), .Y(n1798) );
  AOI22XL U2195 ( .A0(n1761), .A1(y[24]), .B0(n1760), .B1(y[30]), .Y(n1800) );
  AOI221XL U2196 ( .A0(x[67]), .A1(n1968), .B0(x[68]), .B1(n1757), .C0(n1941), 
        .Y(n1942) );
  OAI22XL U2197 ( .A0(x[67]), .A1(n1968), .B0(n1757), .B1(x[68]), .Y(n1941) );
  NOR2XL U2198 ( .A(move_out[2]), .B(n2293), .Y(n2283) );
  NOR2XL U2199 ( .A(move_out[2]), .B(n2286), .Y(n2289) );
  NOR2XL U2200 ( .A(move_out[0]), .B(n2927), .Y(n2288) );
  NOR2XL U2201 ( .A(move_out[1]), .B(n2874), .Y(n2287) );
  NOR2XL U2202 ( .A(move_out[2]), .B(n2295), .Y(n2284) );
  INVXL U2203 ( .A(n2394), .Y(n2393) );
  NAND2XL U2204 ( .A(n2452), .B(n2451), .Y(n2527) );
  NOR2XL U2205 ( .A(n2452), .B(n2451), .Y(n2526) );
  INVXL U2206 ( .A(n2537), .Y(n2525) );
  NOR3XL U2207 ( .A(n2541), .B(n2539), .C(n2531), .Y(n2535) );
  NOR3XL U2208 ( .A(n2542), .B(n2538), .C(n2525), .Y(n2536) );
  INVXL U2209 ( .A(n2543), .Y(n2531) );
  NAND2XL U2210 ( .A(n2511), .B(n2510), .Y(n2519) );
  AOI22XL U2211 ( .A0(n2509), .A1(n2508), .B0(n2507), .B1(n2506), .Y(n2510) );
  AOI22XL U2212 ( .A0(x[73]), .A1(n2497), .B0(n2496), .B1(n2495), .Y(n2511) );
  NAND2XL U2213 ( .A(n2472), .B(n2471), .Y(n2523) );
  AOI22XL U2214 ( .A0(x[74]), .A1(n2497), .B0(n2496), .B1(n2460), .Y(n2472) );
  AOI22XL U2215 ( .A0(n2509), .A1(n2470), .B0(n2507), .B1(n2469), .Y(n2471) );
  AOI21XL U2216 ( .A0(n2507), .A1(n2416), .B0(n2415), .Y(n2517) );
  NAND4XL U2217 ( .A(n2398), .B(n2397), .C(n2396), .D(n2395), .Y(n2416) );
  AOI211XL U2218 ( .A0(n2707), .A1(have_tried_direction[55]), .B0(n2071), .C0(
        n2070), .Y(n2072) );
  NAND2XL U2219 ( .A(n2065), .B(n2064), .Y(n2071) );
  NAND4XL U2220 ( .A(n2069), .B(n2068), .C(n2067), .D(n2066), .Y(n2070) );
  AOI22XL U2221 ( .A0(n2674), .A1(have_tried_direction[199]), .B0(n2755), .B1(
        have_tried_direction[71]), .Y(n2065) );
  AOI22XL U2222 ( .A0(n2181), .A1(have_tried_direction[95]), .B0(n2180), .B1(
        have_tried_direction[119]), .Y(n2061) );
  AOI22XL U2223 ( .A0(n2699), .A1(have_tried_direction[7]), .B0(n2184), .B1(
        have_tried_direction[111]), .Y(n2059) );
  AOI22XL U2224 ( .A0(n2183), .A1(have_tried_direction[79]), .B0(n2182), .B1(
        have_tried_direction[103]), .Y(n2060) );
  AOI22XL U2225 ( .A0(n1768), .A1(have_tried_direction[167]), .B0(n2177), .B1(
        have_tried_direction[175]), .Y(n2074) );
  AOI22XL U2226 ( .A0(n2684), .A1(have_tried_direction[31]), .B0(n2176), .B1(
        have_tried_direction[183]), .Y(n2075) );
  NAND4XL U2227 ( .A(n2204), .B(n2203), .C(n2202), .D(n2201), .Y(n2205) );
  AOI22XL U2228 ( .A0(n2684), .A1(have_tried_direction[24]), .B0(n2176), .B1(
        have_tried_direction[176]), .Y(n2204) );
  AOI22XL U2229 ( .A0(n1768), .A1(have_tried_direction[160]), .B0(n2177), .B1(
        have_tried_direction[168]), .Y(n2203) );
  NAND4XL U2230 ( .A(n2175), .B(n2174), .C(n2173), .D(n2172), .Y(n2206) );
  AOI22XL U2231 ( .A0(n2684), .A1(have_tried_direction[25]), .B0(n2176), .B1(
        have_tried_direction[177]), .Y(n2175) );
  AOI22XL U2232 ( .A0(n1768), .A1(have_tried_direction[161]), .B0(n2177), .B1(
        have_tried_direction[169]), .Y(n2174) );
  NAND4XL U2233 ( .A(n2159), .B(n2158), .C(n2157), .D(n2156), .Y(n2207) );
  AOI22XL U2234 ( .A0(n2684), .A1(have_tried_direction[26]), .B0(n2176), .B1(
        have_tried_direction[178]), .Y(n2159) );
  AOI22XL U2235 ( .A0(n1768), .A1(have_tried_direction[162]), .B0(n2177), .B1(
        have_tried_direction[170]), .Y(n2158) );
  NAND4XL U2236 ( .A(n2143), .B(n2142), .C(n2141), .D(n2140), .Y(n2208) );
  AOI22XL U2237 ( .A0(n2684), .A1(have_tried_direction[27]), .B0(n2176), .B1(
        have_tried_direction[179]), .Y(n2143) );
  AOI22XL U2238 ( .A0(n1768), .A1(have_tried_direction[163]), .B0(n2177), .B1(
        have_tried_direction[171]), .Y(n2142) );
  NAND4XL U2239 ( .A(n2123), .B(n2122), .C(n2121), .D(n2120), .Y(n2124) );
  AOI22XL U2240 ( .A0(n2684), .A1(have_tried_direction[28]), .B0(n2176), .B1(
        have_tried_direction[180]), .Y(n2123) );
  AOI22XL U2241 ( .A0(n1768), .A1(have_tried_direction[164]), .B0(n2177), .B1(
        have_tried_direction[172]), .Y(n2122) );
  NAND4XL U2242 ( .A(n2107), .B(n2106), .C(n2105), .D(n2104), .Y(n2125) );
  AOI22XL U2243 ( .A0(n2684), .A1(have_tried_direction[29]), .B0(n2176), .B1(
        have_tried_direction[181]), .Y(n2107) );
  AOI22XL U2244 ( .A0(n1768), .A1(have_tried_direction[165]), .B0(n2177), .B1(
        have_tried_direction[173]), .Y(n2106) );
  NAND4XL U2245 ( .A(n2091), .B(n2090), .C(n2089), .D(n2088), .Y(n2126) );
  AOI22XL U2246 ( .A0(n2684), .A1(have_tried_direction[30]), .B0(n2176), .B1(
        have_tried_direction[182]), .Y(n2091) );
  AOI22XL U2247 ( .A0(n1768), .A1(have_tried_direction[166]), .B0(n2177), .B1(
        have_tried_direction[174]), .Y(n2090) );
  AOI211XL U2248 ( .A0(n1978), .A1(y[40]), .B0(n1972), .C0(n1971), .Y(n2233)
         );
  AOI22XL U2249 ( .A0(n2892), .A1(n1759), .B0(x[39]), .B1(n1758), .Y(n1967) );
  AOI211XL U2250 ( .A0(n1978), .A1(y[37]), .B0(n1966), .C0(n1965), .Y(n2232)
         );
  AOI22XL U2251 ( .A0(n2901), .A1(n1759), .B0(x[36]), .B1(n1758), .Y(n1962) );
  AOI211XL U2252 ( .A0(n1978), .A1(y[43]), .B0(n1977), .C0(n1976), .Y(n2234)
         );
  AOI22XL U2253 ( .A0(n2902), .A1(n1759), .B0(x[42]), .B1(n1758), .Y(n1973) );
  AOI211XL U2254 ( .A0(n1978), .A1(y[52]), .B0(n1983), .C0(n1982), .Y(n2235)
         );
  AOI22XL U2255 ( .A0(n2888), .A1(n1759), .B0(x[51]), .B1(n1758), .Y(n1979) );
  AOI211XL U2256 ( .A0(y[47]), .A1(n2236), .B0(n2050), .C0(n2049), .Y(n2051)
         );
  NAND4XL U2257 ( .A(n2048), .B(n2047), .C(n2046), .D(n2045), .Y(n2049) );
  AOI22XL U2258 ( .A0(y[50]), .A1(n2237), .B0(y[56]), .B1(n2230), .Y(n2004) );
  AOI211XL U2259 ( .A0(n1978), .A1(y[61]), .B0(n1954), .C0(n1953), .Y(n2256)
         );
  AOI22XL U2260 ( .A0(n2904), .A1(n1759), .B0(x[60]), .B1(n1758), .Y(n1950) );
  AOI211XL U2261 ( .A0(n1978), .A1(y[64]), .B0(n1959), .C0(n1958), .Y(n2257)
         );
  AOI22XL U2262 ( .A0(n2887), .A1(n1759), .B0(x[63]), .B1(n1758), .Y(n1955) );
  OAI21XL U2263 ( .A0(n1978), .A1(y[73]), .B0(n1949), .Y(n2259) );
  AOI211XL U2264 ( .A0(n1978), .A1(y[73]), .B0(n1948), .C0(n1947), .Y(n1949)
         );
  AOI211XL U2265 ( .A0(n1978), .A1(y[1]), .B0(n1889), .C0(n1888), .Y(n2212) );
  AOI22XL U2266 ( .A0(n2883), .A1(n1759), .B0(x[0]), .B1(n1758), .Y(n1829) );
  AOI211XL U2267 ( .A0(n1978), .A1(y[10]), .B0(n1898), .C0(n1897), .Y(n1899)
         );
  OAI21XL U2268 ( .A0(n1978), .A1(y[4]), .B0(n1904), .Y(n2214) );
  AOI211XL U2269 ( .A0(n1978), .A1(y[4]), .B0(n1903), .C0(n1902), .Y(n1904) );
  NOR2XL U2270 ( .A(n2515), .B(n2879), .Y(n1908) );
  NAND2XL U2271 ( .A(n1930), .B(n2518), .Y(n1907) );
  AOI22XL U2272 ( .A0(n1933), .A1(n2878), .B0(direction[2]), .B1(n2518), .Y(
        n1935) );
  NOR2XL U2273 ( .A(n1933), .B(n1929), .Y(n1932) );
  NAND2X1 U2274 ( .A(n1808), .B(n1807), .Y(n1910) );
  AOI22XL U2275 ( .A0(n1916), .A1(y[72]), .B0(n2681), .B1(n1796), .Y(n1808) );
  AOI22XL U2276 ( .A0(n2714), .A1(n1806), .B0(n2721), .B1(n1805), .Y(n1807) );
  NAND4XL U2277 ( .A(n1795), .B(n1794), .C(n1793), .D(n1792), .Y(n1796) );
  NOR2XL U2278 ( .A(direction[1]), .B(n2864), .Y(n2269) );
  NOR2XL U2279 ( .A(direction[0]), .B(n2879), .Y(n2270) );
  AOI211XL U2280 ( .A0(n2801), .A1(in_x[2]), .B0(n2800), .C0(n2799), .Y(n2802)
         );
  NOR2XL U2281 ( .A(n2798), .B(n2797), .Y(n2800) );
  AOI211XL U2282 ( .A0(n2801), .A1(in_y[1]), .B0(n2795), .C0(n2799), .Y(n2796)
         );
  NOR2XL U2283 ( .A(n1978), .B(n2797), .Y(n2795) );
  AOI211XL U2284 ( .A0(n2801), .A1(in_y[0]), .B0(n2686), .C0(n2799), .Y(n2687)
         );
  NOR2XL U2285 ( .A(n2685), .B(n2797), .Y(n2686) );
  AOI211XL U2286 ( .A0(n2801), .A1(in_x[0]), .B0(n2787), .C0(n2799), .Y(n2788)
         );
  NOR2XL U2287 ( .A(n1758), .B(n2797), .Y(n2787) );
  NAND2XL U2288 ( .A(n2808), .B(n2283), .Y(n2775) );
  NAND2XL U2289 ( .A(n2288), .B(n2283), .Y(n2783) );
  NAND2XL U2290 ( .A(n2287), .B(n2283), .Y(n2779) );
  NAND2XL U2291 ( .A(n2289), .B(n2808), .Y(n2767) );
  NAND2XL U2292 ( .A(n2289), .B(n2288), .Y(n2763) );
  NAND2XL U2293 ( .A(n2287), .B(n2289), .Y(n2770) );
  NAND2XL U2294 ( .A(n2288), .B(n2284), .Y(n2757) );
  NAND2XL U2295 ( .A(n2287), .B(n2284), .Y(n2748) );
  AOI211XL U2296 ( .A0(n2801), .A1(in_y[2]), .B0(n2689), .C0(n2799), .Y(n2690)
         );
  NOR2XL U2297 ( .A(n2688), .B(n2797), .Y(n2689) );
  NOR2BXL U2298 ( .AN(n2661), .B(n1595), .Y(n2673) );
  INVX1 U2299 ( .A(n2775), .Y(n2574) );
  INVX1 U2300 ( .A(n2783), .Y(n2575) );
  INVX1 U2301 ( .A(n2779), .Y(n2579) );
  CLKINVX2 U2302 ( .A(n1767), .Y(n2727) );
  NAND2XL U2303 ( .A(direction[1]), .B(direction[0]), .Y(n2573) );
  INVXL U2304 ( .A(n2270), .Y(n2571) );
  INVXL U2305 ( .A(n2269), .Y(n2572) );
  NOR2XL U2306 ( .A(direction[2]), .B(n2573), .Y(n2586) );
  INVXL U2307 ( .A(n2591), .Y(n2585) );
  NAND2XL U2308 ( .A(n2399), .B(n1763), .Y(n2637) );
  NAND2XL U2309 ( .A(n2399), .B(n1762), .Y(n2629) );
  CLKINVX2 U2310 ( .A(n2636), .Y(n2695) );
  NAND2XL U2311 ( .A(n2399), .B(n1767), .Y(n2636) );
  NAND2XL U2312 ( .A(n2399), .B(n1765), .Y(n2634) );
  NAND2XL U2313 ( .A(n2399), .B(n2058), .Y(n2640) );
  INVX1 U2314 ( .A(n2757), .Y(n2630) );
  NAND2XL U2315 ( .A(n1859), .B(n2399), .Y(n2631) );
  CLKINVX2 U2316 ( .A(n2633), .Y(n2750) );
  NAND2XL U2317 ( .A(n2399), .B(n1761), .Y(n2633) );
  NOR3XL U2318 ( .A(direction[1]), .B(direction[0]), .C(n2878), .Y(n2588) );
  NOR2XL U2319 ( .A(direction[2]), .B(n2571), .Y(n2590) );
  NOR2XL U2320 ( .A(direction[2]), .B(n2572), .Y(n2592) );
  INVXL U2321 ( .A(n2526), .Y(n2529) );
  NOR2XL U2322 ( .A(n2526), .B(n2455), .Y(n2532) );
  NAND2XL U2323 ( .A(n2530), .B(n2454), .Y(n2453) );
  AOI31XL U2324 ( .A0(n2536), .A1(n2535), .A2(n2562), .B0(n2534), .Y(n2557) );
  NOR2XL U2325 ( .A(n2547), .B(n2559), .Y(n2534) );
  NAND4XL U2326 ( .A(n2525), .B(n2535), .C(n2542), .D(n2538), .Y(n2556) );
  NAND2XL U2327 ( .A(n2533), .B(n2539), .Y(n2559) );
  NAND2XL U2328 ( .A(n2532), .B(n2531), .Y(n2547) );
  NOR2BXL U2329 ( .AN(n2538), .B(n2537), .Y(n2540) );
  NAND2XL U2330 ( .A(n2543), .B(n2562), .Y(n2558) );
  OAI21XL U2331 ( .A0(n2226), .A1(n2688), .B0(n2225), .Y(n2227) );
  OAI21XL U2332 ( .A0(n2688), .A1(y[71]), .B0(n2224), .Y(n2225) );
  AOI21XL U2333 ( .A0(n1968), .A1(n1758), .B0(n2798), .Y(n2228) );
  NAND4XL U2334 ( .A(n2127), .B(n2126), .C(n2125), .D(n2124), .Y(n2210) );
  NAND4XL U2335 ( .A(n2208), .B(n2207), .C(n2206), .D(n2205), .Y(n2209) );
  NAND4XL U2336 ( .A(n2075), .B(n2074), .C(n2073), .D(n2072), .Y(n2127) );
  NAND3XL U2337 ( .A(n2053), .B(n2052), .C(n2051), .Y(n2054) );
  AOI22XL U2338 ( .A0(y[44]), .A1(n2234), .B0(y[53]), .B1(n2235), .Y(n2052) );
  AOI22XL U2339 ( .A0(y[38]), .A1(n2232), .B0(y[41]), .B1(n2233), .Y(n2053) );
  AOI21XL U2340 ( .A0(y[68]), .A1(n2261), .B0(n1961), .Y(n2056) );
  OAI21XL U2341 ( .A0(n2908), .A1(n2259), .B0(n1960), .Y(n1961) );
  AOI22XL U2342 ( .A0(y[62]), .A1(n2256), .B0(y[65]), .B1(n2257), .Y(n1960) );
  AOI211XL U2343 ( .A0(n2212), .A1(n2913), .B0(n1906), .C0(n1905), .Y(n2057)
         );
  NOR2XL U2344 ( .A(y[8]), .B(n2216), .Y(n1906) );
  OAI22XL U2345 ( .A0(y[11]), .A1(n2211), .B0(y[5]), .B1(n2214), .Y(n1905) );
  OAI21XL U2346 ( .A0(n2264), .A1(n2263), .B0(n2688), .Y(n2265) );
  INVXL U2347 ( .A(n2262), .Y(n2263) );
  NAND2BXL U2348 ( .AN(n2255), .B(n2254), .Y(n2264) );
  AOI22XL U2349 ( .A0(pri[2]), .A1(n2554), .B0(pri[1]), .B1(n2391), .Y(n2271)
         );
  NOR2XL U2350 ( .A(n2270), .B(n2269), .Y(n2391) );
  NOR3XL U2351 ( .A(direction[1]), .B(direction[0]), .C(direction[2]), .Y(
        n2589) );
  AOI211XL U2352 ( .A0(x[53]), .A1(n2579), .B0(n2334), .C0(n2333), .Y(n2335)
         );
  NAND4XL U2353 ( .A(n2332), .B(n2331), .C(n2330), .D(n2329), .Y(n2333) );
  AOI22XL U2354 ( .A0(x[56]), .A1(n2575), .B0(x[59]), .B1(n2574), .Y(n2336) );
  AOI22XL U2355 ( .A0(x[20]), .A1(n2706), .B0(x[17]), .B1(n2694), .Y(n2337) );
  AOI22XL U2356 ( .A0(x[14]), .A1(n2702), .B0(x[23]), .B1(n2710), .Y(n2338) );
  AOI22XL U2357 ( .A0(x[44]), .A1(n2734), .B0(x[41]), .B1(n2737), .Y(n2326) );
  AOI211XL U2358 ( .A0(x[52]), .A1(n2579), .B0(n2350), .C0(n2349), .Y(n2351)
         );
  NAND4XL U2359 ( .A(n2348), .B(n2347), .C(n2346), .D(n2345), .Y(n2349) );
  AOI22XL U2360 ( .A0(x[55]), .A1(n2575), .B0(x[58]), .B1(n2574), .Y(n2352) );
  AOI22XL U2361 ( .A0(x[19]), .A1(n2706), .B0(x[16]), .B1(n2694), .Y(n2353) );
  AOI22XL U2362 ( .A0(x[13]), .A1(n2702), .B0(x[22]), .B1(n2710), .Y(n2354) );
  AOI22XL U2363 ( .A0(x[43]), .A1(n2734), .B0(x[40]), .B1(n2737), .Y(n2342) );
  AOI211XL U2364 ( .A0(y[52]), .A1(n2579), .B0(n2366), .C0(n2365), .Y(n2367)
         );
  NAND4XL U2365 ( .A(n2364), .B(n2363), .C(n2362), .D(n2361), .Y(n2365) );
  AOI22XL U2366 ( .A0(y[55]), .A1(n2575), .B0(y[58]), .B1(n2574), .Y(n2368) );
  AOI22XL U2367 ( .A0(y[19]), .A1(n2706), .B0(y[16]), .B1(n2694), .Y(n2369) );
  AOI22XL U2368 ( .A0(y[13]), .A1(n2702), .B0(y[22]), .B1(n2710), .Y(n2370) );
  AOI22XL U2369 ( .A0(y[43]), .A1(n2734), .B0(y[40]), .B1(n2737), .Y(n2358) );
  AOI211XL U2370 ( .A0(y[51]), .A1(n2579), .B0(n2383), .C0(n2382), .Y(n2384)
         );
  NAND4XL U2371 ( .A(n2381), .B(n2380), .C(n2379), .D(n2378), .Y(n2382) );
  AOI22XL U2372 ( .A0(y[54]), .A1(n2575), .B0(y[57]), .B1(n2574), .Y(n2385) );
  AOI22XL U2373 ( .A0(y[18]), .A1(n2706), .B0(y[15]), .B1(n2694), .Y(n2386) );
  AOI22XL U2374 ( .A0(y[12]), .A1(n2702), .B0(y[21]), .B1(n2710), .Y(n2387) );
  AOI22XL U2375 ( .A0(y[42]), .A1(n2734), .B0(y[39]), .B1(n2737), .Y(n2375) );
  AOI211XL U2376 ( .A0(x[6]), .A1(n2630), .B0(n2318), .C0(n2317), .Y(n2319) );
  NAND4XL U2377 ( .A(n2316), .B(n2315), .C(n2314), .D(n2313), .Y(n2317) );
  AOI22XL U2378 ( .A0(x[54]), .A1(n2575), .B0(x[57]), .B1(n2574), .Y(n2320) );
  AOI22XL U2379 ( .A0(x[18]), .A1(n2706), .B0(x[15]), .B1(n2694), .Y(n2321) );
  AOI22XL U2380 ( .A0(x[12]), .A1(n2702), .B0(x[21]), .B1(n2710), .Y(n2322) );
  AOI22XL U2381 ( .A0(x[42]), .A1(n2734), .B0(x[39]), .B1(n2737), .Y(n2310) );
  AOI211XL U2382 ( .A0(y[53]), .A1(n2579), .B0(n2302), .C0(n2301), .Y(n2303)
         );
  NAND4XL U2383 ( .A(n2300), .B(n2299), .C(n2298), .D(n2297), .Y(n2301) );
  AOI22XL U2384 ( .A0(y[56]), .A1(n2575), .B0(y[59]), .B1(n2574), .Y(n2304) );
  AOI22XL U2385 ( .A0(y[20]), .A1(n2706), .B0(y[17]), .B1(n2694), .Y(n2305) );
  AOI22XL U2386 ( .A0(y[14]), .A1(n2702), .B0(y[23]), .B1(n2710), .Y(n2306) );
  AOI22XL U2387 ( .A0(y[44]), .A1(n2734), .B0(y[41]), .B1(n2737), .Y(n2281) );
  CLKINVX2 U2388 ( .A(n1595), .Y(n2672) );
  NOR2XL U2389 ( .A(n2873), .B(n2292), .Y(n2810) );
  NOR2XL U2390 ( .A(move_out[0]), .B(move_out[1]), .Y(n2807) );
  AOI211XL U2391 ( .A0(n2793), .A1(n1763), .B0(n2792), .C0(n2791), .Y(n2794)
         );
  NOR2XL U2392 ( .A(n2790), .B(n2789), .Y(n2791) );
  AOI31X1 U2393 ( .A0(n2674), .A1(n1766), .A2(n2760), .B0(n2673), .Y(n2806) );
  INVXL U2394 ( .A(n2806), .Y(n2805) );
  CLKINVX2 U2395 ( .A(n2794), .Y(n2837) );
  AOI211XL U2396 ( .A0(n2793), .A1(n1762), .B0(n2723), .C0(n2722), .Y(n2724)
         );
  NOR2XL U2397 ( .A(n2732), .B(n2789), .Y(n2722) );
  INVX1 U2398 ( .A(n2724), .Y(n2836) );
  AOI211XL U2399 ( .A0(n2793), .A1(n2738), .B0(n2726), .C0(n2725), .Y(n2730)
         );
  NOR2XL U2400 ( .A(n2735), .B(n2789), .Y(n2725) );
  INVX1 U2401 ( .A(n2730), .Y(n2835) );
  AOI211XL U2402 ( .A0(n2793), .A1(n1765), .B0(n2729), .C0(n2728), .Y(n2731)
         );
  NOR2XL U2403 ( .A(n2727), .B(n2789), .Y(n2728) );
  INVX1 U2404 ( .A(n2731), .Y(n2834) );
  AOI21XL U2405 ( .A0(n1760), .A1(n2793), .B0(n2777), .Y(n2778) );
  INVX1 U2406 ( .A(n2778), .Y(n2833) );
  AOI21XL U2407 ( .A0(n2785), .A1(n2793), .B0(n2784), .Y(n2786) );
  INVX1 U2408 ( .A(n2786), .Y(n2832) );
  AOI21XL U2409 ( .A0(n1761), .A1(n2793), .B0(n2781), .Y(n2782) );
  INVX1 U2410 ( .A(n2782), .Y(n2831) );
  AOI211XL U2411 ( .A0(n2743), .A1(n2760), .B0(n2742), .C0(n2741), .Y(n2744)
         );
  NOR2XL U2412 ( .A(n2752), .B(n2789), .Y(n2741) );
  INVX1 U2413 ( .A(n2744), .Y(n2830) );
  AOI211XL U2414 ( .A0(n2773), .A1(n1763), .B0(n2746), .C0(n2745), .Y(n2747)
         );
  NOR2XL U2415 ( .A(n2790), .B(n2771), .Y(n2745) );
  INVX1 U2416 ( .A(n2747), .Y(n2829) );
  AOI211XL U2417 ( .A0(n2773), .A1(n1762), .B0(n2734), .C0(n2733), .Y(n2740)
         );
  NOR2XL U2418 ( .A(n2732), .B(n2771), .Y(n2733) );
  INVX1 U2419 ( .A(n2740), .Y(n2828) );
  AOI211XL U2420 ( .A0(n2773), .A1(n2738), .B0(n2737), .C0(n2736), .Y(n2739)
         );
  NOR2XL U2421 ( .A(n2735), .B(n2771), .Y(n2736) );
  INVX1 U2422 ( .A(n2739), .Y(n2827) );
  AOI211XL U2423 ( .A0(n2773), .A1(n1765), .B0(n2716), .C0(n2715), .Y(n2717)
         );
  NOR2XL U2424 ( .A(n2727), .B(n2771), .Y(n2715) );
  INVX1 U2425 ( .A(n2717), .Y(n2826) );
  AOI21XL U2426 ( .A0(n1760), .A1(n2773), .B0(n2768), .Y(n2769) );
  INVX1 U2427 ( .A(n2769), .Y(n2825) );
  AOI21XL U2428 ( .A0(n2765), .A1(n2773), .B0(n2764), .Y(n2766) );
  INVX1 U2429 ( .A(n2766), .Y(n2823) );
  INVX1 U2430 ( .A(n2774), .Y(n2822) );
  AOI211XL U2431 ( .A0(n2755), .A1(n2760), .B0(n2754), .C0(n2753), .Y(n2756)
         );
  NOR2XL U2432 ( .A(n2752), .B(n2771), .Y(n2753) );
  INVX1 U2433 ( .A(n2756), .Y(n2821) );
  AOI211XL U2434 ( .A0(n2711), .A1(n2760), .B0(n2710), .C0(n2709), .Y(n2712)
         );
  NOR2XL U2435 ( .A(n2790), .B(n2758), .Y(n2709) );
  INVX1 U2436 ( .A(n2712), .Y(n2820) );
  AOI211XL U2437 ( .A0(n2707), .A1(n2760), .B0(n2706), .C0(n2705), .Y(n2708)
         );
  NOR2XL U2438 ( .A(n2732), .B(n2758), .Y(n2705) );
  INVX1 U2439 ( .A(n2708), .Y(n2819) );
  AOI211XL U2440 ( .A0(n2695), .A1(n2760), .B0(n2694), .C0(n2693), .Y(n2696)
         );
  NOR2XL U2441 ( .A(n2735), .B(n2758), .Y(n2693) );
  INVX1 U2442 ( .A(n2696), .Y(n2818) );
  AOI211XL U2443 ( .A0(n2703), .A1(n2760), .B0(n2702), .C0(n2701), .Y(n2704)
         );
  NOR2XL U2444 ( .A(n2727), .B(n2758), .Y(n2701) );
  INVX1 U2445 ( .A(n2704), .Y(n2817) );
  AOI21X1 U2446 ( .A0(n2684), .A1(n2760), .B0(n2683), .Y(n2804) );
  INVXL U2447 ( .A(n2804), .Y(n2803) );
  AOI21XL U2448 ( .A0(n2761), .A1(n2760), .B0(n2759), .Y(n2762) );
  INVX1 U2449 ( .A(n2762), .Y(n2816) );
  AOI21XL U2450 ( .A0(n2750), .A1(n2760), .B0(n2749), .Y(n2751) );
  INVX1 U2451 ( .A(n2751), .Y(n2815) );
  AOI211XL U2452 ( .A0(n2699), .A1(n2760), .B0(n2698), .C0(n2697), .Y(n2700)
         );
  NOR2XL U2453 ( .A(n2752), .B(n2758), .Y(n2697) );
  INVX1 U2454 ( .A(n2700), .Y(n2814) );
  NAND2XL U2455 ( .A(n1766), .B(n2674), .Y(n2663) );
  NOR3XL U2456 ( .A(n2573), .B(n2878), .C(n2585), .Y(n2625) );
  NOR3XL U2457 ( .A(n2878), .B(n2571), .C(n2585), .Y(n2622) );
  NOR3XL U2458 ( .A(n2878), .B(n2572), .C(n2585), .Y(n2623) );
  NOR2BXL U2459 ( .AN(n2586), .B(n2585), .Y(n2624) );
  INVXL U2460 ( .A(n2682), .Y(n2639) );
  INVXL U2461 ( .A(n2850), .Y(n2851) );
  INVXL U2462 ( .A(n2855), .Y(n2549) );
  NOR3XL U2463 ( .A(n2873), .B(n2926), .C(n2296), .Y(n2661) );
  NAND2XL U2464 ( .A(n2563), .B(n2850), .Y(n2565) );
  AOI21XL U2465 ( .A0(n2562), .A1(n2561), .B0(n2560), .Y(n2566) );
  INVXL U2466 ( .A(n2556), .Y(n2561) );
  INVXL U2467 ( .A(n2554), .Y(n2555) );
  AND2XL U2468 ( .A(priority_num[2]), .B(n2855), .Y(n2570) );
  INVXL U2469 ( .A(n2532), .Y(n2545) );
  AOI22XL U2470 ( .A0(n2547), .A1(n2558), .B0(n2559), .B1(n2546), .Y(n2563) );
  NAND2XL U2471 ( .A(n2591), .B(n2549), .Y(n2857) );
  NOR2XL U2472 ( .A(n2591), .B(n2855), .Y(n2860) );
  AOI211XL U2473 ( .A0(n2849), .A1(cnt[3]), .B0(n2680), .C0(n2679), .Y(n1597)
         );
  NOR2XL U2474 ( .A(n2678), .B(n2846), .Y(n2679) );
  OAI211XL U2475 ( .A0(move_out[2]), .A1(n2808), .B0(n2672), .C0(n2292), .Y(
        n1603) );
  MXI2XL U2476 ( .A(n2847), .B(n2846), .S0(n2845), .Y(n2848) );
  AOI222XL U2477 ( .A0(n2277), .A1(n2838), .B0(cnt[2]), .B1(n2849), .C0(n2276), 
        .C1(n2720), .Y(n1590) );
  NAND3XL U2478 ( .A(n2578), .B(n1772), .C(n1771), .Y(n2277) );
  AOI211XL U2479 ( .A0(x[50]), .A1(n2742), .B0(n2340), .C0(n2339), .Y(n1580)
         );
  NAND3XL U2480 ( .A(n2327), .B(n2326), .C(n2325), .Y(n2340) );
  NAND4XL U2481 ( .A(n2338), .B(n2337), .C(n2336), .D(n2335), .Y(n2339) );
  AOI22XL U2482 ( .A0(x[26]), .A1(n2754), .B0(x[74]), .B1(n2373), .Y(n2327) );
  AOI211XL U2483 ( .A0(x[49]), .A1(n2742), .B0(n2356), .C0(n2355), .Y(n1581)
         );
  NAND3XL U2484 ( .A(n2343), .B(n2342), .C(n2341), .Y(n2356) );
  NAND4XL U2485 ( .A(n2354), .B(n2353), .C(n2352), .D(n2351), .Y(n2355) );
  AOI211XL U2486 ( .A0(y[49]), .A1(n2742), .B0(n2372), .C0(n2371), .Y(n1582)
         );
  NAND3XL U2487 ( .A(n2359), .B(n2358), .C(n2357), .Y(n2372) );
  NAND4XL U2488 ( .A(n2370), .B(n2369), .C(n2368), .D(n2367), .Y(n2371) );
  AOI211XL U2489 ( .A0(y[48]), .A1(n2742), .B0(n2389), .C0(n2388), .Y(n1583)
         );
  NAND3XL U2490 ( .A(n2376), .B(n2375), .C(n2374), .Y(n2389) );
  NAND4XL U2491 ( .A(n2387), .B(n2386), .C(n2385), .D(n2384), .Y(n2388) );
  AOI211XL U2492 ( .A0(x[48]), .A1(n2742), .B0(n2324), .C0(n2323), .Y(n1584)
         );
  NAND3XL U2493 ( .A(n2311), .B(n2310), .C(n2309), .Y(n2324) );
  NAND4XL U2494 ( .A(n2322), .B(n2321), .C(n2320), .D(n2319), .Y(n2323) );
  AOI211XL U2495 ( .A0(y[50]), .A1(n2742), .B0(n2308), .C0(n2307), .Y(n1586)
         );
  NAND3XL U2496 ( .A(n2282), .B(n2281), .C(n2280), .Y(n2308) );
  NAND4XL U2497 ( .A(n2306), .B(n2305), .C(n2304), .D(n2303), .Y(n2307) );
  AOI2BB2XL U2498 ( .B0(n2824), .B1(n2837), .A0N(n2837), .A1N(x[71]), .Y(n1608) );
  AOI2BB2XL U2499 ( .B0(n2824), .B1(n2836), .A0N(n2836), .A1N(x[68]), .Y(n1611) );
  AOI2BB2XL U2500 ( .B0(n2824), .B1(n2835), .A0N(n2835), .A1N(x[65]), .Y(n1614) );
  AOI2BB2XL U2501 ( .B0(n2824), .B1(n2834), .A0N(n2834), .A1N(x[62]), .Y(n1617) );
  AOI2BB2XL U2502 ( .B0(n2824), .B1(n2833), .A0N(n2833), .A1N(x[59]), .Y(n1620) );
  AOI2BB2XL U2503 ( .B0(n2824), .B1(n2832), .A0N(n2832), .A1N(x[56]), .Y(n1623) );
  AOI2BB2XL U2504 ( .B0(n2824), .B1(n2831), .A0N(n2831), .A1N(x[53]), .Y(n1626) );
  AOI2BB2XL U2505 ( .B0(n2824), .B1(n2830), .A0N(n2830), .A1N(x[50]), .Y(n1629) );
  AOI2BB2XL U2506 ( .B0(n2824), .B1(n2829), .A0N(n2829), .A1N(x[47]), .Y(n1632) );
  AOI2BB2XL U2507 ( .B0(n2824), .B1(n2828), .A0N(n2828), .A1N(x[44]), .Y(n1635) );
  AOI2BB2XL U2508 ( .B0(n2824), .B1(n2827), .A0N(n2827), .A1N(x[41]), .Y(n1638) );
  AOI2BB2XL U2509 ( .B0(n2824), .B1(n2826), .A0N(n2826), .A1N(x[38]), .Y(n1641) );
  AOI2BB2XL U2510 ( .B0(n2824), .B1(n2825), .A0N(n2825), .A1N(x[35]), .Y(n1644) );
  AOI2BB2XL U2511 ( .B0(n2824), .B1(n2823), .A0N(n2823), .A1N(x[32]), .Y(n1647) );
  AOI2BB2XL U2512 ( .B0(n2824), .B1(n2822), .A0N(n2822), .A1N(x[29]), .Y(n1650) );
  AOI2BB2XL U2513 ( .B0(n2824), .B1(n2821), .A0N(n2821), .A1N(x[26]), .Y(n1653) );
  AOI2BB2XL U2514 ( .B0(n2824), .B1(n2820), .A0N(n2820), .A1N(x[23]), .Y(n1656) );
  AOI2BB2XL U2515 ( .B0(n2824), .B1(n2819), .A0N(n2819), .A1N(x[20]), .Y(n1659) );
  AOI2BB2XL U2516 ( .B0(n2824), .B1(n2818), .A0N(n2818), .A1N(x[17]), .Y(n1662) );
  AOI2BB2XL U2517 ( .B0(n2824), .B1(n2817), .A0N(n2817), .A1N(x[14]), .Y(n1665) );
  AOI22XL U2518 ( .A0(n2804), .A1(n2930), .B0(n2824), .B1(n2803), .Y(n1668) );
  AOI2BB2XL U2519 ( .B0(n2824), .B1(n2816), .A0N(n2816), .A1N(x[8]), .Y(n1671)
         );
  AOI2BB2XL U2520 ( .B0(n2824), .B1(n2815), .A0N(n2815), .A1N(x[5]), .Y(n1674)
         );
  AOI2BB2XL U2521 ( .B0(n2824), .B1(n2814), .A0N(n2814), .A1N(x[2]), .Y(n1677)
         );
  AOI22XL U2522 ( .A0(n2806), .A1(n2880), .B0(n2824), .B1(n2805), .Y(n1755) );
  AOI22XL U2523 ( .A0(n2806), .A1(n2877), .B0(n2813), .B1(n2805), .Y(n1606) );
  AOI2BB2XL U2524 ( .B0(n2813), .B1(n2837), .A0N(n2837), .A1N(x[70]), .Y(n1609) );
  AOI2BB2XL U2525 ( .B0(n2813), .B1(n2836), .A0N(n2836), .A1N(x[67]), .Y(n1612) );
  AOI2BB2XL U2526 ( .B0(n2813), .B1(n2835), .A0N(n2835), .A1N(x[64]), .Y(n1615) );
  AOI2BB2XL U2527 ( .B0(n2813), .B1(n2834), .A0N(n2834), .A1N(x[61]), .Y(n1618) );
  AOI2BB2XL U2528 ( .B0(n2813), .B1(n2833), .A0N(n2833), .A1N(x[58]), .Y(n1621) );
  AOI2BB2XL U2529 ( .B0(n2813), .B1(n2832), .A0N(n2832), .A1N(x[55]), .Y(n1624) );
  AOI2BB2XL U2530 ( .B0(n2813), .B1(n2831), .A0N(n2831), .A1N(x[52]), .Y(n1627) );
  AOI2BB2XL U2531 ( .B0(n2813), .B1(n2830), .A0N(n2830), .A1N(x[49]), .Y(n1630) );
  AOI2BB2XL U2532 ( .B0(n2813), .B1(n2829), .A0N(n2829), .A1N(x[46]), .Y(n1633) );
  AOI2BB2XL U2533 ( .B0(n2813), .B1(n2828), .A0N(n2828), .A1N(x[43]), .Y(n1636) );
  AOI2BB2XL U2534 ( .B0(n2813), .B1(n2827), .A0N(n2827), .A1N(x[40]), .Y(n1639) );
  AOI2BB2XL U2535 ( .B0(n2813), .B1(n2826), .A0N(n2826), .A1N(x[37]), .Y(n1642) );
  AOI2BB2XL U2536 ( .B0(n2813), .B1(n2825), .A0N(n2825), .A1N(x[34]), .Y(n1645) );
  AOI2BB2XL U2537 ( .B0(n2813), .B1(n2823), .A0N(n2823), .A1N(x[31]), .Y(n1648) );
  AOI2BB2XL U2538 ( .B0(n2813), .B1(n2822), .A0N(n2822), .A1N(x[28]), .Y(n1651) );
  AOI2BB2XL U2539 ( .B0(n2813), .B1(n2821), .A0N(n2821), .A1N(x[25]), .Y(n1654) );
  AOI2BB2XL U2540 ( .B0(n2813), .B1(n2820), .A0N(n2820), .A1N(x[22]), .Y(n1657) );
  AOI2BB2XL U2541 ( .B0(n2813), .B1(n2819), .A0N(n2819), .A1N(x[19]), .Y(n1660) );
  AOI2BB2XL U2542 ( .B0(n2813), .B1(n2818), .A0N(n2818), .A1N(x[16]), .Y(n1663) );
  AOI2BB2XL U2543 ( .B0(n2813), .B1(n2817), .A0N(n2817), .A1N(x[13]), .Y(n1666) );
  AOI22XL U2544 ( .A0(n2804), .A1(n2931), .B0(n2813), .B1(n2803), .Y(n1669) );
  AOI2BB2XL U2545 ( .B0(n2813), .B1(n2816), .A0N(n2816), .A1N(x[7]), .Y(n1672)
         );
  AOI2BB2XL U2546 ( .B0(n2813), .B1(n2815), .A0N(n2815), .A1N(x[4]), .Y(n1675)
         );
  AOI2BB2XL U2547 ( .B0(n2813), .B1(n2814), .A0N(n2814), .A1N(x[1]), .Y(n1678)
         );
  AOI22XL U2548 ( .A0(n2806), .A1(n2910), .B0(n2811), .B1(n2805), .Y(n1681) );
  AOI2BB2XL U2549 ( .B0(n2811), .B1(n2837), .A0N(n2837), .A1N(y[70]), .Y(n1684) );
  AOI2BB2XL U2550 ( .B0(n2811), .B1(n2836), .A0N(n2836), .A1N(y[67]), .Y(n1687) );
  AOI2BB2XL U2551 ( .B0(n2811), .B1(n2835), .A0N(n2835), .A1N(y[64]), .Y(n1690) );
  AOI2BB2XL U2552 ( .B0(n2811), .B1(n2834), .A0N(n2834), .A1N(y[61]), .Y(n1693) );
  AOI2BB2XL U2553 ( .B0(n2811), .B1(n2833), .A0N(n2833), .A1N(y[58]), .Y(n1696) );
  AOI2BB2XL U2554 ( .B0(n2811), .B1(n2832), .A0N(n2832), .A1N(y[55]), .Y(n1699) );
  AOI2BB2XL U2555 ( .B0(n2811), .B1(n2831), .A0N(n2831), .A1N(y[52]), .Y(n1702) );
  AOI2BB2XL U2556 ( .B0(n2811), .B1(n2830), .A0N(n2830), .A1N(y[49]), .Y(n1705) );
  AOI2BB2XL U2557 ( .B0(n2811), .B1(n2829), .A0N(n2829), .A1N(y[46]), .Y(n1708) );
  AOI2BB2XL U2558 ( .B0(n2811), .B1(n2828), .A0N(n2828), .A1N(y[43]), .Y(n1711) );
  AOI2BB2XL U2559 ( .B0(n2811), .B1(n2827), .A0N(n2827), .A1N(y[40]), .Y(n1714) );
  AOI2BB2XL U2560 ( .B0(n2811), .B1(n2826), .A0N(n2826), .A1N(y[37]), .Y(n1717) );
  AOI2BB2XL U2561 ( .B0(n2811), .B1(n2825), .A0N(n2825), .A1N(y[34]), .Y(n1720) );
  AOI2BB2XL U2562 ( .B0(n2811), .B1(n2823), .A0N(n2823), .A1N(y[31]), .Y(n1723) );
  AOI2BB2XL U2563 ( .B0(n2811), .B1(n2822), .A0N(n2822), .A1N(y[28]), .Y(n1726) );
  AOI2BB2XL U2564 ( .B0(n2811), .B1(n2821), .A0N(n2821), .A1N(y[25]), .Y(n1729) );
  AOI2BB2XL U2565 ( .B0(n2811), .B1(n2820), .A0N(n2820), .A1N(y[22]), .Y(n1732) );
  AOI2BB2XL U2566 ( .B0(n2811), .B1(n2819), .A0N(n2819), .A1N(y[19]), .Y(n1735) );
  AOI2BB2XL U2567 ( .B0(n2811), .B1(n2818), .A0N(n2818), .A1N(y[16]), .Y(n1738) );
  AOI2BB2XL U2568 ( .B0(n2811), .B1(n2817), .A0N(n2817), .A1N(y[13]), .Y(n1741) );
  AOI22XL U2569 ( .A0(n2804), .A1(n2928), .B0(n2811), .B1(n2803), .Y(n1744) );
  AOI2BB2XL U2570 ( .B0(n2811), .B1(n2816), .A0N(n2816), .A1N(y[7]), .Y(n1747)
         );
  AOI2BB2XL U2571 ( .B0(n2811), .B1(n2815), .A0N(n2815), .A1N(y[4]), .Y(n1750)
         );
  AOI2BB2XL U2572 ( .B0(n2811), .B1(n2814), .A0N(n2814), .A1N(y[1]), .Y(n1753)
         );
  AOI22XL U2573 ( .A0(n2806), .A1(n2886), .B0(n2692), .B1(n2805), .Y(n1682) );
  AOI2BB2XL U2574 ( .B0(n2692), .B1(n2837), .A0N(n2837), .A1N(y[69]), .Y(n1685) );
  AOI22XL U2575 ( .A0(n2724), .A1(n2895), .B0(n2692), .B1(n2836), .Y(n1688) );
  AOI22XL U2576 ( .A0(n2730), .A1(n2887), .B0(n2692), .B1(n2835), .Y(n1691) );
  AOI22XL U2577 ( .A0(n2731), .A1(n2904), .B0(n2692), .B1(n2834), .Y(n1694) );
  AOI22XL U2578 ( .A0(n2778), .A1(n2893), .B0(n2692), .B1(n2833), .Y(n1697) );
  AOI22XL U2579 ( .A0(n2786), .A1(n2903), .B0(n2692), .B1(n2832), .Y(n1700) );
  AOI22XL U2580 ( .A0(n2782), .A1(n2888), .B0(n2692), .B1(n2831), .Y(n1703) );
  AOI22XL U2581 ( .A0(n2744), .A1(n2882), .B0(n2692), .B1(n2830), .Y(n1706) );
  AOI22XL U2582 ( .A0(n2747), .A1(n2885), .B0(n2692), .B1(n2829), .Y(n1709) );
  AOI22XL U2583 ( .A0(n2740), .A1(n2902), .B0(n2692), .B1(n2828), .Y(n1712) );
  AOI22XL U2584 ( .A0(n2739), .A1(n2892), .B0(n2692), .B1(n2827), .Y(n1715) );
  AOI22XL U2585 ( .A0(n2717), .A1(n2901), .B0(n2692), .B1(n2826), .Y(n1718) );
  AOI22XL U2586 ( .A0(n2769), .A1(n2891), .B0(n2692), .B1(n2825), .Y(n1721) );
  AOI22XL U2587 ( .A0(n2766), .A1(n2900), .B0(n2692), .B1(n2823), .Y(n1724) );
  AOI22XL U2588 ( .A0(n2774), .A1(n2896), .B0(n2692), .B1(n2822), .Y(n1727) );
  AOI22XL U2589 ( .A0(n2756), .A1(n2889), .B0(n2692), .B1(n2821), .Y(n1730) );
  AOI22XL U2590 ( .A0(n2712), .A1(n2884), .B0(n2692), .B1(n2820), .Y(n1733) );
  AOI22XL U2591 ( .A0(n2708), .A1(n2899), .B0(n2692), .B1(n2819), .Y(n1736) );
  AOI22XL U2592 ( .A0(n2696), .A1(n2890), .B0(n2692), .B1(n2818), .Y(n1739) );
  AOI22XL U2593 ( .A0(n2704), .A1(n2898), .B0(n2692), .B1(n2817), .Y(n1742) );
  AOI22XL U2594 ( .A0(n2804), .A1(n2881), .B0(n2692), .B1(n2803), .Y(n1745) );
  AOI22XL U2595 ( .A0(n2762), .A1(n2897), .B0(n2692), .B1(n2816), .Y(n1748) );
  AOI22XL U2596 ( .A0(n2751), .A1(n2894), .B0(n2692), .B1(n2815), .Y(n1751) );
  AOI22XL U2597 ( .A0(n2700), .A1(n2883), .B0(n2692), .B1(n2814), .Y(n1754) );
  AOI22XL U2598 ( .A0(n2806), .A1(n2911), .B0(n2812), .B1(n2805), .Y(n1607) );
  AOI22XL U2599 ( .A0(n2794), .A1(n2905), .B0(n2812), .B1(n2837), .Y(n1610) );
  AOI2BB2XL U2600 ( .B0(n2812), .B1(n2836), .A0N(n2836), .A1N(x[66]), .Y(n1613) );
  AOI2BB2XL U2601 ( .B0(n2812), .B1(n2835), .A0N(n2835), .A1N(x[63]), .Y(n1616) );
  AOI2BB2XL U2602 ( .B0(n2812), .B1(n2834), .A0N(n2834), .A1N(x[60]), .Y(n1619) );
  AOI2BB2XL U2603 ( .B0(n2812), .B1(n2833), .A0N(n2833), .A1N(x[57]), .Y(n1622) );
  AOI2BB2XL U2604 ( .B0(n2812), .B1(n2832), .A0N(n2832), .A1N(x[54]), .Y(n1625) );
  AOI2BB2XL U2605 ( .B0(n2812), .B1(n2831), .A0N(n2831), .A1N(x[51]), .Y(n1628) );
  AOI2BB2XL U2606 ( .B0(n2812), .B1(n2830), .A0N(n2830), .A1N(x[48]), .Y(n1631) );
  AOI2BB2XL U2607 ( .B0(n2812), .B1(n2829), .A0N(n2829), .A1N(x[45]), .Y(n1634) );
  AOI2BB2XL U2608 ( .B0(n2812), .B1(n2828), .A0N(n2828), .A1N(x[42]), .Y(n1637) );
  AOI2BB2XL U2609 ( .B0(n2812), .B1(n2827), .A0N(n2827), .A1N(x[39]), .Y(n1640) );
  AOI2BB2XL U2610 ( .B0(n2812), .B1(n2826), .A0N(n2826), .A1N(x[36]), .Y(n1643) );
  AOI2BB2XL U2611 ( .B0(n2812), .B1(n2825), .A0N(n2825), .A1N(x[33]), .Y(n1646) );
  AOI2BB2XL U2612 ( .B0(n2812), .B1(n2823), .A0N(n2823), .A1N(x[30]), .Y(n1649) );
  AOI2BB2XL U2613 ( .B0(n2812), .B1(n2822), .A0N(n2822), .A1N(x[27]), .Y(n1652) );
  AOI2BB2XL U2614 ( .B0(n2812), .B1(n2821), .A0N(n2821), .A1N(x[24]), .Y(n1655) );
  AOI2BB2XL U2615 ( .B0(n2812), .B1(n2820), .A0N(n2820), .A1N(x[21]), .Y(n1658) );
  AOI2BB2XL U2616 ( .B0(n2812), .B1(n2819), .A0N(n2819), .A1N(x[18]), .Y(n1661) );
  AOI2BB2XL U2617 ( .B0(n2812), .B1(n2818), .A0N(n2818), .A1N(x[15]), .Y(n1664) );
  AOI2BB2XL U2618 ( .B0(n2812), .B1(n2817), .A0N(n2817), .A1N(x[12]), .Y(n1667) );
  AOI22XL U2619 ( .A0(n2804), .A1(n2929), .B0(n2812), .B1(n2803), .Y(n1670) );
  AOI2BB2XL U2620 ( .B0(n2812), .B1(n2816), .A0N(n2816), .A1N(x[6]), .Y(n1673)
         );
  AOI2BB2XL U2621 ( .B0(n2812), .B1(n2815), .A0N(n2815), .A1N(x[3]), .Y(n1676)
         );
  AOI2BB2XL U2622 ( .B0(n2812), .B1(n2814), .A0N(n2814), .A1N(x[0]), .Y(n1679)
         );
  AOI22XL U2623 ( .A0(n2806), .A1(n2908), .B0(n2691), .B1(n2805), .Y(n1680) );
  AOI2BB2XL U2624 ( .B0(n2691), .B1(n2837), .A0N(n2837), .A1N(y[71]), .Y(n1683) );
  AOI22XL U2625 ( .A0(n2724), .A1(n2915), .B0(n2691), .B1(n2836), .Y(n1686) );
  AOI22XL U2626 ( .A0(n2730), .A1(n2872), .B0(n2691), .B1(n2835), .Y(n1689) );
  AOI22XL U2627 ( .A0(n2731), .A1(n2922), .B0(n2691), .B1(n2834), .Y(n1692) );
  AOI22XL U2628 ( .A0(n2778), .A1(n2909), .B0(n2691), .B1(n2833), .Y(n1695) );
  AOI22XL U2629 ( .A0(n2786), .A1(n2907), .B0(n2691), .B1(n2832), .Y(n1698) );
  AOI22XL U2630 ( .A0(n2782), .A1(n2867), .B0(n2691), .B1(n2831), .Y(n1701) );
  AOI22XL U2631 ( .A0(n2744), .A1(n2865), .B0(n2691), .B1(n2830), .Y(n1704) );
  AOI22XL U2632 ( .A0(n2747), .A1(n2914), .B0(n2691), .B1(n2829), .Y(n1707) );
  AOI22XL U2633 ( .A0(n2740), .A1(n2921), .B0(n2691), .B1(n2828), .Y(n1710) );
  AOI22XL U2634 ( .A0(n2739), .A1(n2871), .B0(n2691), .B1(n2827), .Y(n1713) );
  AOI22XL U2635 ( .A0(n2717), .A1(n2920), .B0(n2691), .B1(n2826), .Y(n1716) );
  AOI22XL U2636 ( .A0(n2769), .A1(n2870), .B0(n2691), .B1(n2825), .Y(n1719) );
  AOI22XL U2637 ( .A0(n2766), .A1(n2868), .B0(n2691), .B1(n2823), .Y(n1722) );
  AOI22XL U2638 ( .A0(n2774), .A1(n2917), .B0(n2691), .B1(n2822), .Y(n1725) );
  AOI22XL U2639 ( .A0(n2756), .A1(n2916), .B0(n2691), .B1(n2821), .Y(n1728) );
  AOI22XL U2640 ( .A0(n2712), .A1(n2866), .B0(n2691), .B1(n2820), .Y(n1731) );
  AOI22XL U2641 ( .A0(n2708), .A1(n2919), .B0(n2691), .B1(n2819), .Y(n1734) );
  AOI22XL U2642 ( .A0(n2696), .A1(n2869), .B0(n2691), .B1(n2818), .Y(n1737) );
  AOI22XL U2643 ( .A0(n2704), .A1(n2918), .B0(n2691), .B1(n2817), .Y(n1740) );
  AOI22XL U2644 ( .A0(n2804), .A1(n2906), .B0(n2691), .B1(n2803), .Y(n1743) );
  AOI22XL U2645 ( .A0(n2762), .A1(n2923), .B0(n2691), .B1(n2816), .Y(n1746) );
  AOI22XL U2646 ( .A0(n2751), .A1(n2912), .B0(n2691), .B1(n2815), .Y(n1749) );
  AOI22XL U2647 ( .A0(n2700), .A1(n2913), .B0(n2691), .B1(n2814), .Y(n1752) );
  AOI22XL U2648 ( .A0(have_tried_direction[199]), .A1(n2669), .B0(n2584), .B1(
        n2667), .Y(n1381) );
  AOI22XL U2649 ( .A0(have_tried_direction[198]), .A1(n2669), .B0(n2577), .B1(
        n2667), .Y(n1382) );
  AOI22XL U2650 ( .A0(have_tried_direction[197]), .A1(n2669), .B0(n2583), .B1(
        n2667), .Y(n1383) );
  AOI22XL U2651 ( .A0(have_tried_direction[196]), .A1(n2669), .B0(n2664), .B1(
        n2667), .Y(n1384) );
  AOI22XL U2652 ( .A0(have_tried_direction[195]), .A1(n2669), .B0(n2587), .B1(
        n2667), .Y(n1385) );
  AOI22XL U2653 ( .A0(have_tried_direction[194]), .A1(n2669), .B0(n2668), .B1(
        n2667), .Y(n1386) );
  AOI22XL U2654 ( .A0(have_tried_direction[193]), .A1(n2669), .B0(n2666), .B1(
        n2667), .Y(n1387) );
  AOI22XL U2655 ( .A0(have_tried_direction[192]), .A1(n2669), .B0(n2665), .B1(
        n2667), .Y(n1388) );
  AOI22XL U2656 ( .A0(have_tried_direction[191]), .A1(n2616), .B0(n2584), .B1(
        n2615), .Y(n1389) );
  AOI22XL U2657 ( .A0(have_tried_direction[190]), .A1(n2616), .B0(n2577), .B1(
        n2615), .Y(n1390) );
  AOI22XL U2658 ( .A0(have_tried_direction[189]), .A1(n2616), .B0(n2583), .B1(
        n2615), .Y(n1391) );
  AOI22XL U2659 ( .A0(have_tried_direction[188]), .A1(n2616), .B0(n2664), .B1(
        n2615), .Y(n1392) );
  AOI22XL U2660 ( .A0(have_tried_direction[187]), .A1(n2616), .B0(n2587), .B1(
        n2615), .Y(n1393) );
  AOI22XL U2661 ( .A0(have_tried_direction[186]), .A1(n2616), .B0(n2668), .B1(
        n2615), .Y(n1394) );
  AOI22XL U2662 ( .A0(have_tried_direction[185]), .A1(n2616), .B0(n2666), .B1(
        n2615), .Y(n1395) );
  AOI22XL U2663 ( .A0(have_tried_direction[184]), .A1(n2616), .B0(n2665), .B1(
        n2615), .Y(n1396) );
  AOI22XL U2664 ( .A0(have_tried_direction[183]), .A1(n2618), .B0(n2584), .B1(
        n2617), .Y(n1397) );
  AOI22XL U2665 ( .A0(have_tried_direction[182]), .A1(n2618), .B0(n2577), .B1(
        n2617), .Y(n1398) );
  AOI22XL U2666 ( .A0(have_tried_direction[181]), .A1(n2618), .B0(n2583), .B1(
        n2617), .Y(n1399) );
  AOI22XL U2667 ( .A0(have_tried_direction[180]), .A1(n2618), .B0(n2664), .B1(
        n2617), .Y(n1400) );
  AOI22XL U2668 ( .A0(have_tried_direction[179]), .A1(n2618), .B0(n2587), .B1(
        n2617), .Y(n1401) );
  AOI22XL U2669 ( .A0(have_tried_direction[178]), .A1(n2618), .B0(n2668), .B1(
        n2617), .Y(n1402) );
  AOI22XL U2670 ( .A0(have_tried_direction[177]), .A1(n2618), .B0(n2666), .B1(
        n2617), .Y(n1403) );
  AOI22XL U2671 ( .A0(have_tried_direction[176]), .A1(n2618), .B0(n2665), .B1(
        n2617), .Y(n1404) );
  AOI22XL U2672 ( .A0(have_tried_direction[175]), .A1(n2614), .B0(n2584), .B1(
        n2613), .Y(n1405) );
  AOI22XL U2673 ( .A0(have_tried_direction[174]), .A1(n2614), .B0(n2577), .B1(
        n2613), .Y(n1406) );
  AOI22XL U2674 ( .A0(have_tried_direction[173]), .A1(n2614), .B0(n2583), .B1(
        n2613), .Y(n1407) );
  AOI22XL U2675 ( .A0(have_tried_direction[172]), .A1(n2614), .B0(n2664), .B1(
        n2613), .Y(n1408) );
  AOI22XL U2676 ( .A0(have_tried_direction[171]), .A1(n2614), .B0(n2587), .B1(
        n2613), .Y(n1409) );
  AOI22XL U2677 ( .A0(have_tried_direction[170]), .A1(n2614), .B0(n2668), .B1(
        n2613), .Y(n1410) );
  AOI22XL U2678 ( .A0(have_tried_direction[169]), .A1(n2614), .B0(n2666), .B1(
        n2613), .Y(n1411) );
  AOI22XL U2679 ( .A0(have_tried_direction[168]), .A1(n2614), .B0(n2665), .B1(
        n2613), .Y(n1412) );
  AOI22XL U2680 ( .A0(have_tried_direction[167]), .A1(n2608), .B0(n2584), .B1(
        n2607), .Y(n1413) );
  AOI22XL U2681 ( .A0(have_tried_direction[166]), .A1(n2608), .B0(n2577), .B1(
        n2607), .Y(n1414) );
  AOI22XL U2682 ( .A0(have_tried_direction[165]), .A1(n2608), .B0(n2583), .B1(
        n2607), .Y(n1415) );
  AOI22XL U2683 ( .A0(have_tried_direction[164]), .A1(n2608), .B0(n2664), .B1(
        n2607), .Y(n1416) );
  AOI22XL U2684 ( .A0(have_tried_direction[163]), .A1(n2608), .B0(n2587), .B1(
        n2607), .Y(n1417) );
  AOI22XL U2685 ( .A0(have_tried_direction[162]), .A1(n2608), .B0(n2668), .B1(
        n2607), .Y(n1418) );
  AOI22XL U2686 ( .A0(have_tried_direction[161]), .A1(n2608), .B0(n2666), .B1(
        n2607), .Y(n1419) );
  AOI22XL U2687 ( .A0(have_tried_direction[160]), .A1(n2608), .B0(n2665), .B1(
        n2607), .Y(n1420) );
  AOI22XL U2688 ( .A0(have_tried_direction[159]), .A1(n2602), .B0(n2584), .B1(
        n2601), .Y(n1421) );
  AOI22XL U2689 ( .A0(have_tried_direction[158]), .A1(n2602), .B0(n2577), .B1(
        n2601), .Y(n1422) );
  AOI22XL U2690 ( .A0(have_tried_direction[157]), .A1(n2602), .B0(n2583), .B1(
        n2601), .Y(n1423) );
  AOI22XL U2691 ( .A0(have_tried_direction[156]), .A1(n2602), .B0(n2664), .B1(
        n2601), .Y(n1424) );
  AOI22XL U2692 ( .A0(have_tried_direction[155]), .A1(n2602), .B0(n2587), .B1(
        n2601), .Y(n1425) );
  AOI22XL U2693 ( .A0(have_tried_direction[154]), .A1(n2602), .B0(n2668), .B1(
        n2601), .Y(n1426) );
  AOI22XL U2694 ( .A0(have_tried_direction[153]), .A1(n2602), .B0(n2666), .B1(
        n2601), .Y(n1427) );
  AOI22XL U2695 ( .A0(have_tried_direction[152]), .A1(n2602), .B0(n2665), .B1(
        n2601), .Y(n1428) );
  AOI22XL U2696 ( .A0(have_tried_direction[151]), .A1(n2610), .B0(n2584), .B1(
        n2609), .Y(n1429) );
  AOI22XL U2697 ( .A0(have_tried_direction[150]), .A1(n2610), .B0(n2577), .B1(
        n2609), .Y(n1430) );
  AOI22XL U2698 ( .A0(have_tried_direction[149]), .A1(n2610), .B0(n2583), .B1(
        n2609), .Y(n1431) );
  AOI22XL U2699 ( .A0(have_tried_direction[148]), .A1(n2610), .B0(n2664), .B1(
        n2609), .Y(n1432) );
  AOI22XL U2700 ( .A0(have_tried_direction[147]), .A1(n2610), .B0(n2587), .B1(
        n2609), .Y(n1433) );
  AOI22XL U2701 ( .A0(have_tried_direction[146]), .A1(n2610), .B0(n2668), .B1(
        n2609), .Y(n1434) );
  AOI22XL U2702 ( .A0(have_tried_direction[145]), .A1(n2610), .B0(n2666), .B1(
        n2609), .Y(n1435) );
  AOI22XL U2703 ( .A0(have_tried_direction[144]), .A1(n2610), .B0(n2665), .B1(
        n2609), .Y(n1436) );
  AOI22XL U2704 ( .A0(have_tried_direction[143]), .A1(n2606), .B0(n2584), .B1(
        n2605), .Y(n1437) );
  AOI22XL U2705 ( .A0(have_tried_direction[142]), .A1(n2606), .B0(n2577), .B1(
        n2605), .Y(n1438) );
  AOI22XL U2706 ( .A0(have_tried_direction[141]), .A1(n2606), .B0(n2583), .B1(
        n2605), .Y(n1439) );
  AOI22XL U2707 ( .A0(have_tried_direction[140]), .A1(n2606), .B0(n2664), .B1(
        n2605), .Y(n1440) );
  AOI22XL U2708 ( .A0(have_tried_direction[139]), .A1(n2606), .B0(n2587), .B1(
        n2605), .Y(n1441) );
  AOI22XL U2709 ( .A0(have_tried_direction[138]), .A1(n2606), .B0(n2668), .B1(
        n2605), .Y(n1442) );
  AOI22XL U2710 ( .A0(have_tried_direction[137]), .A1(n2606), .B0(n2666), .B1(
        n2605), .Y(n1443) );
  AOI22XL U2711 ( .A0(have_tried_direction[136]), .A1(n2606), .B0(n2665), .B1(
        n2605), .Y(n1444) );
  AOI22XL U2712 ( .A0(have_tried_direction[135]), .A1(n2648), .B0(n2584), .B1(
        n2647), .Y(n1445) );
  AOI22XL U2713 ( .A0(have_tried_direction[134]), .A1(n2648), .B0(n2577), .B1(
        n2647), .Y(n1446) );
  AOI22XL U2714 ( .A0(have_tried_direction[133]), .A1(n2648), .B0(n2583), .B1(
        n2647), .Y(n1447) );
  AOI22XL U2715 ( .A0(have_tried_direction[132]), .A1(n2648), .B0(n2664), .B1(
        n2647), .Y(n1448) );
  AOI22XL U2716 ( .A0(have_tried_direction[131]), .A1(n2648), .B0(n2587), .B1(
        n2647), .Y(n1449) );
  AOI22XL U2717 ( .A0(have_tried_direction[130]), .A1(n2648), .B0(n2668), .B1(
        n2647), .Y(n1450) );
  AOI22XL U2718 ( .A0(have_tried_direction[129]), .A1(n2648), .B0(n2666), .B1(
        n2647), .Y(n1451) );
  AOI22XL U2719 ( .A0(have_tried_direction[128]), .A1(n2648), .B0(n2665), .B1(
        n2647), .Y(n1452) );
  AOI22XL U2720 ( .A0(have_tried_direction[127]), .A1(n2612), .B0(n2584), .B1(
        n2611), .Y(n1453) );
  AOI22XL U2721 ( .A0(have_tried_direction[126]), .A1(n2612), .B0(n2577), .B1(
        n2611), .Y(n1454) );
  AOI22XL U2722 ( .A0(have_tried_direction[125]), .A1(n2612), .B0(n2583), .B1(
        n2611), .Y(n1455) );
  AOI22XL U2723 ( .A0(have_tried_direction[124]), .A1(n2612), .B0(n2664), .B1(
        n2611), .Y(n1456) );
  AOI22XL U2724 ( .A0(have_tried_direction[123]), .A1(n2612), .B0(n2587), .B1(
        n2611), .Y(n1457) );
  AOI22XL U2725 ( .A0(have_tried_direction[122]), .A1(n2612), .B0(n2668), .B1(
        n2611), .Y(n1458) );
  AOI22XL U2726 ( .A0(have_tried_direction[121]), .A1(n2612), .B0(n2666), .B1(
        n2611), .Y(n1459) );
  AOI22XL U2727 ( .A0(have_tried_direction[120]), .A1(n2612), .B0(n2665), .B1(
        n2611), .Y(n1460) );
  AOI22XL U2728 ( .A0(have_tried_direction[119]), .A1(n2604), .B0(n2584), .B1(
        n2603), .Y(n1461) );
  AOI22XL U2729 ( .A0(have_tried_direction[118]), .A1(n2604), .B0(n2577), .B1(
        n2603), .Y(n1462) );
  AOI22XL U2730 ( .A0(have_tried_direction[117]), .A1(n2604), .B0(n2583), .B1(
        n2603), .Y(n1463) );
  AOI22XL U2731 ( .A0(have_tried_direction[116]), .A1(n2604), .B0(n2664), .B1(
        n2603), .Y(n1464) );
  AOI22XL U2732 ( .A0(have_tried_direction[115]), .A1(n2604), .B0(n2587), .B1(
        n2603), .Y(n1465) );
  AOI22XL U2733 ( .A0(have_tried_direction[114]), .A1(n2604), .B0(n2668), .B1(
        n2603), .Y(n1466) );
  AOI22XL U2734 ( .A0(have_tried_direction[113]), .A1(n2604), .B0(n2666), .B1(
        n2603), .Y(n1467) );
  AOI22XL U2735 ( .A0(have_tried_direction[112]), .A1(n2604), .B0(n2665), .B1(
        n2603), .Y(n1468) );
  AOI22XL U2736 ( .A0(have_tried_direction[111]), .A1(n2600), .B0(n2584), .B1(
        n2599), .Y(n1469) );
  AOI22XL U2737 ( .A0(have_tried_direction[110]), .A1(n2600), .B0(n2577), .B1(
        n2599), .Y(n1470) );
  AOI22XL U2738 ( .A0(have_tried_direction[109]), .A1(n2600), .B0(n2583), .B1(
        n2599), .Y(n1471) );
  AOI22XL U2739 ( .A0(have_tried_direction[108]), .A1(n2600), .B0(n2664), .B1(
        n2599), .Y(n1472) );
  AOI22XL U2740 ( .A0(have_tried_direction[107]), .A1(n2600), .B0(n2587), .B1(
        n2599), .Y(n1473) );
  AOI22XL U2741 ( .A0(have_tried_direction[106]), .A1(n2600), .B0(n2668), .B1(
        n2599), .Y(n1474) );
  AOI22XL U2742 ( .A0(have_tried_direction[105]), .A1(n2600), .B0(n2666), .B1(
        n2599), .Y(n1475) );
  AOI22XL U2743 ( .A0(have_tried_direction[104]), .A1(n2600), .B0(n2665), .B1(
        n2599), .Y(n1476) );
  AOI22XL U2744 ( .A0(have_tried_direction[103]), .A1(n2594), .B0(n2584), .B1(
        n2593), .Y(n1477) );
  AOI22XL U2745 ( .A0(have_tried_direction[102]), .A1(n2594), .B0(n2577), .B1(
        n2593), .Y(n1478) );
  AOI22XL U2746 ( .A0(have_tried_direction[101]), .A1(n2594), .B0(n2583), .B1(
        n2593), .Y(n1479) );
  AOI22XL U2747 ( .A0(have_tried_direction[100]), .A1(n2594), .B0(n2664), .B1(
        n2593), .Y(n1480) );
  AOI22XL U2748 ( .A0(have_tried_direction[99]), .A1(n2594), .B0(n2587), .B1(
        n2593), .Y(n1481) );
  AOI22XL U2749 ( .A0(have_tried_direction[98]), .A1(n2594), .B0(n2668), .B1(
        n2593), .Y(n1482) );
  AOI22XL U2750 ( .A0(have_tried_direction[97]), .A1(n2594), .B0(n2666), .B1(
        n2593), .Y(n1483) );
  AOI22XL U2751 ( .A0(have_tried_direction[96]), .A1(n2594), .B0(n2665), .B1(
        n2593), .Y(n1484) );
  AOI22XL U2752 ( .A0(have_tried_direction[95]), .A1(n2596), .B0(n2584), .B1(
        n2595), .Y(n1485) );
  AOI22XL U2753 ( .A0(have_tried_direction[94]), .A1(n2596), .B0(n2577), .B1(
        n2595), .Y(n1486) );
  AOI22XL U2754 ( .A0(have_tried_direction[93]), .A1(n2596), .B0(n2583), .B1(
        n2595), .Y(n1487) );
  AOI22XL U2755 ( .A0(have_tried_direction[92]), .A1(n2596), .B0(n2664), .B1(
        n2595), .Y(n1488) );
  AOI22XL U2756 ( .A0(have_tried_direction[91]), .A1(n2596), .B0(n2587), .B1(
        n2595), .Y(n1489) );
  AOI22XL U2757 ( .A0(have_tried_direction[90]), .A1(n2596), .B0(n2668), .B1(
        n2595), .Y(n1490) );
  AOI22XL U2758 ( .A0(have_tried_direction[89]), .A1(n2596), .B0(n2666), .B1(
        n2595), .Y(n1491) );
  AOI22XL U2759 ( .A0(have_tried_direction[88]), .A1(n2596), .B0(n2665), .B1(
        n2595), .Y(n1492) );
  AOI22XL U2760 ( .A0(have_tried_direction[87]), .A1(n2598), .B0(n2584), .B1(
        n2597), .Y(n1493) );
  AOI22XL U2761 ( .A0(have_tried_direction[86]), .A1(n2598), .B0(n2577), .B1(
        n2597), .Y(n1494) );
  AOI22XL U2762 ( .A0(have_tried_direction[85]), .A1(n2598), .B0(n2583), .B1(
        n2597), .Y(n1495) );
  AOI22XL U2763 ( .A0(have_tried_direction[84]), .A1(n2598), .B0(n2664), .B1(
        n2597), .Y(n1496) );
  AOI22XL U2764 ( .A0(have_tried_direction[83]), .A1(n2598), .B0(n2587), .B1(
        n2597), .Y(n1497) );
  AOI22XL U2765 ( .A0(have_tried_direction[82]), .A1(n2598), .B0(n2668), .B1(
        n2597), .Y(n1498) );
  AOI22XL U2766 ( .A0(have_tried_direction[81]), .A1(n2598), .B0(n2666), .B1(
        n2597), .Y(n1499) );
  AOI22XL U2767 ( .A0(have_tried_direction[80]), .A1(n2598), .B0(n2665), .B1(
        n2597), .Y(n1500) );
  AOI22XL U2768 ( .A0(have_tried_direction[79]), .A1(n2627), .B0(n2626), .B1(
        n2625), .Y(n1501) );
  AOI22XL U2769 ( .A0(have_tried_direction[78]), .A1(n2627), .B0(n2626), .B1(
        n2622), .Y(n1502) );
  AOI22XL U2770 ( .A0(have_tried_direction[77]), .A1(n2627), .B0(n2626), .B1(
        n2623), .Y(n1503) );
  AOI22XL U2771 ( .A0(have_tried_direction[76]), .A1(n2627), .B0(n2626), .B1(
        n2664), .Y(n1504) );
  AOI22XL U2772 ( .A0(have_tried_direction[75]), .A1(n2627), .B0(n2626), .B1(
        n2624), .Y(n1505) );
  AOI22XL U2773 ( .A0(have_tried_direction[74]), .A1(n2627), .B0(n2626), .B1(
        n2668), .Y(n1506) );
  AOI22XL U2774 ( .A0(have_tried_direction[73]), .A1(n2627), .B0(n2626), .B1(
        n2666), .Y(n1507) );
  AOI22XL U2775 ( .A0(have_tried_direction[72]), .A1(n2627), .B0(n2665), .B1(
        n2626), .Y(n1508) );
  AOI22XL U2776 ( .A0(have_tried_direction[71]), .A1(n2658), .B0(n2584), .B1(
        n2657), .Y(n1509) );
  AOI22XL U2777 ( .A0(have_tried_direction[70]), .A1(n2658), .B0(n2577), .B1(
        n2657), .Y(n1510) );
  AOI22XL U2778 ( .A0(have_tried_direction[69]), .A1(n2658), .B0(n2583), .B1(
        n2657), .Y(n1511) );
  AOI22XL U2779 ( .A0(have_tried_direction[68]), .A1(n2658), .B0(n2664), .B1(
        n2657), .Y(n1512) );
  AOI22XL U2780 ( .A0(have_tried_direction[67]), .A1(n2658), .B0(n2587), .B1(
        n2657), .Y(n1513) );
  AOI22XL U2781 ( .A0(have_tried_direction[66]), .A1(n2658), .B0(n2668), .B1(
        n2657), .Y(n1514) );
  AOI22XL U2782 ( .A0(have_tried_direction[65]), .A1(n2658), .B0(n2666), .B1(
        n2657), .Y(n1515) );
  AOI22XL U2783 ( .A0(have_tried_direction[64]), .A1(n2658), .B0(n2665), .B1(
        n2657), .Y(n1516) );
  AOI22XL U2784 ( .A0(have_tried_direction[63]), .A1(n2654), .B0(n2584), .B1(
        n2653), .Y(n1517) );
  AOI22XL U2785 ( .A0(have_tried_direction[62]), .A1(n2654), .B0(n2577), .B1(
        n2653), .Y(n1518) );
  AOI22XL U2786 ( .A0(have_tried_direction[61]), .A1(n2654), .B0(n2583), .B1(
        n2653), .Y(n1519) );
  AOI22XL U2787 ( .A0(have_tried_direction[60]), .A1(n2654), .B0(n2664), .B1(
        n2653), .Y(n1520) );
  AOI22XL U2788 ( .A0(have_tried_direction[59]), .A1(n2654), .B0(n2587), .B1(
        n2653), .Y(n1521) );
  AOI22XL U2789 ( .A0(have_tried_direction[58]), .A1(n2654), .B0(n2668), .B1(
        n2653), .Y(n1522) );
  AOI22XL U2790 ( .A0(have_tried_direction[57]), .A1(n2654), .B0(n2666), .B1(
        n2653), .Y(n1523) );
  AOI22XL U2791 ( .A0(have_tried_direction[56]), .A1(n2654), .B0(n2665), .B1(
        n2653), .Y(n1524) );
  AOI22XL U2792 ( .A0(have_tried_direction[55]), .A1(n2656), .B0(n2584), .B1(
        n2655), .Y(n1525) );
  AOI22XL U2793 ( .A0(have_tried_direction[54]), .A1(n2656), .B0(n2577), .B1(
        n2655), .Y(n1526) );
  AOI22XL U2794 ( .A0(have_tried_direction[53]), .A1(n2656), .B0(n2583), .B1(
        n2655), .Y(n1527) );
  AOI22XL U2795 ( .A0(have_tried_direction[52]), .A1(n2656), .B0(n2664), .B1(
        n2655), .Y(n1528) );
  AOI22XL U2796 ( .A0(have_tried_direction[51]), .A1(n2656), .B0(n2587), .B1(
        n2655), .Y(n1529) );
  AOI22XL U2797 ( .A0(have_tried_direction[50]), .A1(n2656), .B0(n2668), .B1(
        n2655), .Y(n1530) );
  AOI22XL U2798 ( .A0(have_tried_direction[49]), .A1(n2656), .B0(n2666), .B1(
        n2655), .Y(n1531) );
  AOI22XL U2799 ( .A0(have_tried_direction[48]), .A1(n2656), .B0(n2665), .B1(
        n2655), .Y(n1532) );
  AOI22XL U2800 ( .A0(have_tried_direction[47]), .A1(n2646), .B0(n2584), .B1(
        n2645), .Y(n1533) );
  AOI22XL U2801 ( .A0(have_tried_direction[46]), .A1(n2646), .B0(n2577), .B1(
        n2645), .Y(n1534) );
  AOI22XL U2802 ( .A0(have_tried_direction[45]), .A1(n2646), .B0(n2583), .B1(
        n2645), .Y(n1535) );
  AOI22XL U2803 ( .A0(have_tried_direction[44]), .A1(n2646), .B0(n2664), .B1(
        n2645), .Y(n1536) );
  AOI22XL U2804 ( .A0(have_tried_direction[43]), .A1(n2646), .B0(n2587), .B1(
        n2645), .Y(n1537) );
  AOI22XL U2805 ( .A0(have_tried_direction[42]), .A1(n2646), .B0(n2668), .B1(
        n2645), .Y(n1538) );
  AOI22XL U2806 ( .A0(have_tried_direction[41]), .A1(n2646), .B0(n2666), .B1(
        n2645), .Y(n1539) );
  AOI22XL U2807 ( .A0(have_tried_direction[40]), .A1(n2646), .B0(n2665), .B1(
        n2645), .Y(n1540) );
  AOI22XL U2808 ( .A0(have_tried_direction[39]), .A1(n2650), .B0(n2584), .B1(
        n2649), .Y(n1541) );
  AOI22XL U2809 ( .A0(have_tried_direction[38]), .A1(n2650), .B0(n2577), .B1(
        n2649), .Y(n1542) );
  AOI22XL U2810 ( .A0(have_tried_direction[37]), .A1(n2650), .B0(n2583), .B1(
        n2649), .Y(n1543) );
  AOI22XL U2811 ( .A0(have_tried_direction[36]), .A1(n2650), .B0(n2664), .B1(
        n2649), .Y(n1544) );
  AOI22XL U2812 ( .A0(have_tried_direction[35]), .A1(n2650), .B0(n2587), .B1(
        n2649), .Y(n1545) );
  AOI22XL U2813 ( .A0(have_tried_direction[34]), .A1(n2650), .B0(n2668), .B1(
        n2649), .Y(n1546) );
  AOI22XL U2814 ( .A0(have_tried_direction[33]), .A1(n2650), .B0(n2666), .B1(
        n2649), .Y(n1547) );
  AOI22XL U2815 ( .A0(have_tried_direction[32]), .A1(n2650), .B0(n2665), .B1(
        n2649), .Y(n1548) );
  AOI22XL U2816 ( .A0(have_tried_direction[31]), .A1(n2660), .B0(n2584), .B1(
        n2659), .Y(n1549) );
  AOI22XL U2817 ( .A0(have_tried_direction[30]), .A1(n2660), .B0(n2577), .B1(
        n2659), .Y(n1550) );
  AOI22XL U2818 ( .A0(have_tried_direction[29]), .A1(n2660), .B0(n2583), .B1(
        n2659), .Y(n1551) );
  AOI22XL U2819 ( .A0(have_tried_direction[28]), .A1(n2660), .B0(n2664), .B1(
        n2659), .Y(n1552) );
  AOI22XL U2820 ( .A0(have_tried_direction[27]), .A1(n2660), .B0(n2587), .B1(
        n2659), .Y(n1553) );
  AOI22XL U2821 ( .A0(have_tried_direction[26]), .A1(n2660), .B0(n2668), .B1(
        n2659), .Y(n1554) );
  AOI22XL U2822 ( .A0(have_tried_direction[25]), .A1(n2660), .B0(n2666), .B1(
        n2659), .Y(n1555) );
  AOI22XL U2823 ( .A0(have_tried_direction[24]), .A1(n2660), .B0(n2665), .B1(
        n2659), .Y(n1556) );
  AOI22XL U2824 ( .A0(have_tried_direction[23]), .A1(n2652), .B0(n2584), .B1(
        n2651), .Y(n1557) );
  AOI22XL U2825 ( .A0(have_tried_direction[22]), .A1(n2652), .B0(n2577), .B1(
        n2651), .Y(n1558) );
  AOI22XL U2826 ( .A0(have_tried_direction[21]), .A1(n2652), .B0(n2583), .B1(
        n2651), .Y(n1559) );
  AOI22XL U2827 ( .A0(have_tried_direction[20]), .A1(n2652), .B0(n2664), .B1(
        n2651), .Y(n1560) );
  AOI22XL U2828 ( .A0(have_tried_direction[19]), .A1(n2652), .B0(n2587), .B1(
        n2651), .Y(n1561) );
  AOI22XL U2829 ( .A0(have_tried_direction[18]), .A1(n2652), .B0(n2668), .B1(
        n2651), .Y(n1562) );
  AOI22XL U2830 ( .A0(have_tried_direction[17]), .A1(n2652), .B0(n2666), .B1(
        n2651), .Y(n1563) );
  AOI22XL U2831 ( .A0(have_tried_direction[16]), .A1(n2652), .B0(n2665), .B1(
        n2651), .Y(n1564) );
  AOI22XL U2832 ( .A0(have_tried_direction[15]), .A1(n2644), .B0(n2584), .B1(
        n2643), .Y(n1565) );
  AOI22XL U2833 ( .A0(have_tried_direction[14]), .A1(n2644), .B0(n2577), .B1(
        n2643), .Y(n1566) );
  AOI22XL U2834 ( .A0(have_tried_direction[13]), .A1(n2644), .B0(n2583), .B1(
        n2643), .Y(n1567) );
  AOI22XL U2835 ( .A0(have_tried_direction[12]), .A1(n2644), .B0(n2664), .B1(
        n2643), .Y(n1568) );
  AOI22XL U2836 ( .A0(have_tried_direction[11]), .A1(n2644), .B0(n2587), .B1(
        n2643), .Y(n1569) );
  AOI22XL U2837 ( .A0(have_tried_direction[10]), .A1(n2644), .B0(n2668), .B1(
        n2643), .Y(n1570) );
  AOI22XL U2838 ( .A0(have_tried_direction[9]), .A1(n2644), .B0(n2666), .B1(
        n2643), .Y(n1571) );
  AOI22XL U2839 ( .A0(have_tried_direction[8]), .A1(n2644), .B0(n2665), .B1(
        n2643), .Y(n1572) );
  AOI22XL U2840 ( .A0(have_tried_direction[7]), .A1(n2642), .B0(n2584), .B1(
        n2641), .Y(n1573) );
  AOI22XL U2841 ( .A0(have_tried_direction[6]), .A1(n2642), .B0(n2577), .B1(
        n2641), .Y(n1574) );
  AOI22XL U2842 ( .A0(have_tried_direction[5]), .A1(n2642), .B0(n2583), .B1(
        n2641), .Y(n1575) );
  AOI22XL U2843 ( .A0(have_tried_direction[4]), .A1(n2642), .B0(n2664), .B1(
        n2641), .Y(n1576) );
  AOI22XL U2844 ( .A0(have_tried_direction[3]), .A1(n2642), .B0(n2587), .B1(
        n2641), .Y(n1577) );
  AOI22XL U2845 ( .A0(have_tried_direction[2]), .A1(n2642), .B0(n2668), .B1(
        n2641), .Y(n1578) );
  AOI22XL U2846 ( .A0(have_tried_direction[1]), .A1(n2642), .B0(n2666), .B1(
        n2641), .Y(n1579) );
  NAND2XL U2847 ( .A(n2855), .B(priority_num[0]), .Y(n2856) );
  AOI22XL U2848 ( .A0(n2855), .A1(priority_num[0]), .B0(pri[0]), .B1(n2549), 
        .Y(n1589) );
  AOI31XL U2849 ( .A0(cnt[4]), .A1(n2183), .A2(n2591), .B0(n1770), .Y(n1596)
         );
  OAI22XL U2850 ( .A0(cs[1]), .A1(n2671), .B0(n2661), .B1(n1595), .Y(n1770) );
  AOI211XL U2851 ( .A0(n2860), .A1(direction[2]), .B0(n2570), .C0(n2569), .Y(
        n1598) );
  AOI21XL U2852 ( .A0(n2568), .A1(n2567), .B0(n2857), .Y(n2569) );
  AOI22XL U2853 ( .A0(n2853), .A1(pri[2]), .B0(n2854), .B1(n2555), .Y(n2568)
         );
  AOI211XL U2854 ( .A0(direction[1]), .A1(n2860), .B0(n2553), .C0(n2552), .Y(
        n1599) );
  AOI21XL U2855 ( .A0(n2551), .A1(n2550), .B0(n2857), .Y(n2553) );
  AOI22XL U2856 ( .A0(n2853), .A1(pri[1]), .B0(n2854), .B1(n2392), .Y(n2551)
         );
  AOI22XL U2857 ( .A0(have_tried_direction[0]), .A1(n2642), .B0(n2665), .B1(
        n2641), .Y(n1600) );
  AOI21XL U2858 ( .A0(n2507), .A1(n2450), .B0(n2449), .Y(n2451) );
  NAND2BX4 U2859 ( .AN(n2718), .B(n2638), .Y(n2581) );
  OR3XL U2860 ( .A(n2808), .B(n2807), .C(n1595), .Y(n1604) );
  NOR2X2 U2861 ( .A(n2874), .B(n2927), .Y(n2808) );
  NAND3X2 U2862 ( .A(n2672), .B(n2873), .C(n2926), .Y(n2295) );
  NOR2X2 U2863 ( .A(n2861), .B(n2578), .Y(n2181) );
  CLKINVX3 U2864 ( .A(n2058), .Y(n2578) );
  NAND2BX4 U2865 ( .AN(n2713), .B(n2638), .Y(n2621) );
  NAND2X2 U2866 ( .A(n2862), .B(cnt[3]), .Y(n2713) );
  NOR2X1 U2867 ( .A(n2401), .B(n2400), .Y(n2496) );
  OAI21XL U2868 ( .A0(n2393), .A1(cnt[3]), .B0(cnt[4]), .Y(n2401) );
  NAND2X1 U2869 ( .A(n1595), .B(n2846), .Y(n2799) );
  NOR3X2 U2870 ( .A(n1595), .B(n2873), .C(n2926), .Y(n2373) );
  NAND2X2 U2871 ( .A(cs[0]), .B(cs[1]), .Y(n1595) );
  NOR2X2 U2872 ( .A(n2780), .B(n2862), .Y(n2194) );
  NAND2X2 U2873 ( .A(cnt[4]), .B(n2861), .Y(n2718) );
  NOR2X2 U2874 ( .A(n2861), .B(n2776), .Y(n2182) );
  NOR2X2 U2875 ( .A(n2780), .B(n2861), .Y(n2179) );
  NOR2X4 U2876 ( .A(cnt[1]), .B(n1772), .Y(n1854) );
  AOI21XL U2877 ( .A0(direction[1]), .A1(n2521), .B0(n1848), .Y(n1849) );
  OR3XL U2878 ( .A(cnt[1]), .B(n2875), .C(n2863), .Y(n2063) );
  AOI21XL U2879 ( .A0(n2524), .A1(n1880), .B0(n1879), .Y(n1881) );
  AOI21XL U2880 ( .A0(n2688), .A1(y[71]), .B0(n2223), .Y(n2224) );
  AOI21XL U2881 ( .A0(n2530), .A1(n2529), .B0(n2528), .Y(n2562) );
  AOI21XL U2882 ( .A0(n1761), .A1(n2773), .B0(n2772), .Y(n2774) );
  INVX1 U2883 ( .A(in_valid), .Y(n2671) );
  NOR2X2 U2884 ( .A(cnt[1]), .B(cnt[2]), .Y(n2394) );
  OR2X2 U2885 ( .A(n2863), .B(n2393), .Y(n2752) );
  NOR2X2 U2886 ( .A(n2861), .B(n2752), .Y(n2183) );
  NAND2BX2 U2887 ( .AN(move_out[2]), .B(n2807), .Y(n2296) );
  NAND2X4 U2888 ( .A(n2394), .B(n2863), .Y(n2790) );
  NOR2X2 U2889 ( .A(cnt[3]), .B(cnt[4]), .Y(n2399) );
  NOR2X1 U2890 ( .A(n2635), .B(n2671), .Y(n2855) );
  AOI21XL U2891 ( .A0(pri[1]), .A1(n2549), .B0(n2552), .Y(n1587) );
  AOI21XL U2892 ( .A0(pri[2]), .A1(n2549), .B0(n2570), .Y(n1588) );
  NAND2X1 U2893 ( .A(cnt[2]), .B(n2863), .Y(n1772) );
  NAND2XL U2894 ( .A(cnt[2]), .B(n2876), .Y(n1771) );
  NOR3X2 U2895 ( .A(cnt[2]), .B(N2025), .C(n2876), .Y(n2785) );
  CLKINVX3 U2896 ( .A(n2785), .Y(n2780) );
  OR2X2 U2897 ( .A(n2875), .B(n2844), .Y(n2732) );
  OR2X2 U2898 ( .A(n2876), .B(n1772), .Y(n2735) );
  NOR2X2 U2899 ( .A(n1783), .B(n2842), .Y(n2721) );
  AOI21XL U2900 ( .A0(direction[2]), .A1(n2270), .B0(n2586), .Y(n1930) );
  MX2X1 U2901 ( .A(n2879), .B(direction[1]), .S0(n1910), .Y(n2685) );
  MX2X1 U2902 ( .A(n2879), .B(direction[1]), .S0(n2512), .Y(n2219) );
  OAI221XL U2903 ( .A0(n2883), .A1(n1759), .B0(n1758), .B1(x[0]), .C0(n1829), 
        .Y(n1889) );
  AOI21XL U2904 ( .A0(direction[2]), .A1(n2269), .B0(n2589), .Y(n1873) );
  AOI21X1 U2905 ( .A0(n2714), .A1(n1869), .B0(n1868), .Y(n2524) );
  OAI21XL U2906 ( .A0(n1875), .A1(n1878), .B0(n1874), .Y(n1876) );
  OAI21XL U2907 ( .A0(n1877), .A1(n2512), .B0(n1876), .Y(n1882) );
  OAI21XL U2908 ( .A0(n2524), .A1(n1880), .B0(direction[1]), .Y(n1879) );
  OAI21XL U2909 ( .A0(n1978), .A1(y[1]), .B0(n1887), .Y(n1888) );
  OAI221XL U2910 ( .A0(x[8]), .A1(n1757), .B0(x[7]), .B1(n1968), .C0(n1890), 
        .Y(n1893) );
  OAI221XL U2911 ( .A0(n2897), .A1(n1759), .B0(n1758), .B1(x[6]), .C0(n1891), 
        .Y(n1892) );
  OAI221XL U2912 ( .A0(x[11]), .A1(n1757), .B0(x[10]), .B1(n1968), .C0(n1895), 
        .Y(n1898) );
  OAI221XL U2913 ( .A0(n2881), .A1(n1759), .B0(n1758), .B1(x[9]), .C0(n1896), 
        .Y(n1897) );
  OAI21XL U2914 ( .A0(n1978), .A1(y[10]), .B0(n1899), .Y(n2211) );
  OAI221XL U2915 ( .A0(x[5]), .A1(n1757), .B0(x[4]), .B1(n1968), .C0(n1900), 
        .Y(n1903) );
  OAI221XL U2916 ( .A0(n2894), .A1(n1759), .B0(n1758), .B1(x[3]), .C0(n1901), 
        .Y(n1902) );
  OAI21XL U2917 ( .A0(n1908), .A1(n2518), .B0(n1907), .Y(n1909) );
  CLKINVX3 U2918 ( .A(n2780), .Y(n2765) );
  NAND2X2 U2919 ( .A(n1928), .B(n1927), .Y(n2530) );
  OAI21XL U2920 ( .A0(n2518), .A1(n1930), .B0(n2515), .Y(n1931) );
  OAI21XL U2921 ( .A0(n1932), .A1(n2515), .B0(n1931), .Y(n1937) );
  AOI21XL U2922 ( .A0(n1935), .A1(n2530), .B0(direction[1]), .Y(n1934) );
  OAI21XL U2923 ( .A0(n1935), .A1(n2530), .B0(n1934), .Y(n1936) );
  AOI21X2 U2924 ( .A0(n1939), .A1(n2530), .B0(n1938), .Y(n2688) );
  OAI221XL U2925 ( .A0(n2895), .A1(n1759), .B0(n1758), .B1(x[66]), .C0(n1940), 
        .Y(n1944) );
  OAI21XL U2926 ( .A0(n1978), .A1(y[67]), .B0(n1942), .Y(n1943) );
  OAI221XL U2927 ( .A0(x[73]), .A1(n1968), .B0(n1764), .B1(n2880), .C0(n1945), 
        .Y(n1948) );
  OAI221XL U2928 ( .A0(n2886), .A1(n1759), .B0(n1758), .B1(x[72]), .C0(n1946), 
        .Y(n1947) );
  OAI221XL U2929 ( .A0(n2904), .A1(n1759), .B0(n1758), .B1(x[60]), .C0(n1950), 
        .Y(n1954) );
  OAI21XL U2930 ( .A0(n1978), .A1(y[61]), .B0(n1952), .Y(n1953) );
  OAI221XL U2931 ( .A0(n2887), .A1(n1759), .B0(n1758), .B1(x[63]), .C0(n1955), 
        .Y(n1959) );
  OAI21XL U2932 ( .A0(n1978), .A1(y[64]), .B0(n1957), .Y(n1958) );
  OAI221XL U2933 ( .A0(n2901), .A1(n1759), .B0(n1758), .B1(x[36]), .C0(n1962), 
        .Y(n1966) );
  OAI21XL U2934 ( .A0(n1978), .A1(y[37]), .B0(n1964), .Y(n1965) );
  OAI221XL U2935 ( .A0(n2892), .A1(n1759), .B0(n1758), .B1(x[39]), .C0(n1967), 
        .Y(n1972) );
  OAI21XL U2936 ( .A0(n1978), .A1(y[40]), .B0(n1970), .Y(n1971) );
  OAI221XL U2937 ( .A0(n2902), .A1(n1759), .B0(n1758), .B1(x[42]), .C0(n1973), 
        .Y(n1977) );
  OAI21XL U2938 ( .A0(n1978), .A1(y[43]), .B0(n1975), .Y(n1976) );
  OAI221XL U2939 ( .A0(n2888), .A1(n1759), .B0(n1758), .B1(x[51]), .C0(n1979), 
        .Y(n1983) );
  OAI21XL U2940 ( .A0(n1978), .A1(y[52]), .B0(n1981), .Y(n1982) );
  OAI221XL U2941 ( .A0(n2885), .A1(n1759), .B0(n1758), .B1(x[45]), .C0(n1984), 
        .Y(n1988) );
  OAI21XL U2942 ( .A0(n1978), .A1(y[46]), .B0(n1986), .Y(n1987) );
  OAI221XL U2943 ( .A0(x[59]), .A1(n1757), .B0(x[58]), .B1(n1968), .C0(n1989), 
        .Y(n1992) );
  OAI221XL U2944 ( .A0(n2893), .A1(n1759), .B0(n1758), .B1(x[57]), .C0(n1990), 
        .Y(n1991) );
  OAI21XL U2945 ( .A0(n1978), .A1(y[58]), .B0(n1993), .Y(n2231) );
  OAI221XL U2946 ( .A0(n2882), .A1(n1759), .B0(n1758), .B1(x[48]), .C0(n1994), 
        .Y(n1998) );
  OAI21XL U2947 ( .A0(n1978), .A1(y[49]), .B0(n1996), .Y(n1997) );
  OAI221XL U2948 ( .A0(n2903), .A1(n1759), .B0(n1758), .B1(x[54]), .C0(n1999), 
        .Y(n2003) );
  OAI21XL U2949 ( .A0(n1978), .A1(y[55]), .B0(n2001), .Y(n2002) );
  OAI21XL U2950 ( .A0(n2909), .A1(n2231), .B0(n2004), .Y(n2050) );
  OAI221XL U2951 ( .A0(n2898), .A1(n1759), .B0(n1758), .B1(x[12]), .C0(n2005), 
        .Y(n2009) );
  OAI21XL U2952 ( .A0(n1978), .A1(y[13]), .B0(n2007), .Y(n2008) );
  OAI221XL U2953 ( .A0(n2890), .A1(n1759), .B0(n1758), .B1(x[15]), .C0(n2010), 
        .Y(n2014) );
  OAI21XL U2954 ( .A0(n1978), .A1(y[16]), .B0(n2012), .Y(n2013) );
  OAI221XL U2955 ( .A0(n2899), .A1(n1759), .B0(n1758), .B1(x[18]), .C0(n2015), 
        .Y(n2019) );
  OAI21XL U2956 ( .A0(n1978), .A1(y[19]), .B0(n2017), .Y(n2018) );
  OAI221XL U2957 ( .A0(n2884), .A1(n1759), .B0(n1758), .B1(x[21]), .C0(n2020), 
        .Y(n2024) );
  OAI21XL U2958 ( .A0(n1978), .A1(y[22]), .B0(n2022), .Y(n2023) );
  OAI221XL U2959 ( .A0(n2889), .A1(n1759), .B0(n1758), .B1(x[24]), .C0(n2025), 
        .Y(n2029) );
  OAI21XL U2960 ( .A0(n1978), .A1(y[25]), .B0(n2027), .Y(n2028) );
  OAI221XL U2961 ( .A0(n2900), .A1(n1759), .B0(n1758), .B1(x[30]), .C0(n2030), 
        .Y(n2034) );
  OAI21XL U2962 ( .A0(n1978), .A1(y[31]), .B0(n2032), .Y(n2033) );
  OAI221XL U2963 ( .A0(n2896), .A1(n1759), .B0(n1758), .B1(x[27]), .C0(n2035), 
        .Y(n2039) );
  OAI21XL U2964 ( .A0(n1978), .A1(y[28]), .B0(n2037), .Y(n2038) );
  OAI221XL U2965 ( .A0(n2891), .A1(n1759), .B0(n1758), .B1(x[33]), .C0(n2040), 
        .Y(n2044) );
  OAI21XL U2966 ( .A0(n1978), .A1(y[34]), .B0(n2042), .Y(n2043) );
  AOI21XL U2967 ( .A0(n2685), .A1(n1978), .B0(n2688), .Y(n2229) );
  NOR2X2 U2968 ( .A(n2862), .B(n2735), .Y(n2176) );
  NOR2X2 U2969 ( .A(n2862), .B(n2063), .Y(n2177) );
  NOR2X2 U2970 ( .A(n2861), .B(n2735), .Y(n2180) );
  NOR2X2 U2971 ( .A(n2861), .B(n2063), .Y(n2184) );
  NOR2X2 U2972 ( .A(n2862), .B(n2732), .Y(n2191) );
  NOR2X2 U2973 ( .A(n2861), .B(n2732), .Y(n2840) );
  OAI221XL U2974 ( .A0(x[71]), .A1(n1757), .B0(y[70]), .B1(n1978), .C0(n2217), 
        .Y(n2221) );
  OAI221XL U2975 ( .A0(x[70]), .A1(n1968), .B0(n2905), .B1(n2219), .C0(n2218), 
        .Y(n2220) );
  OAI21XL U2976 ( .A0(y[69]), .A1(n2685), .B0(n2222), .Y(n2223) );
  NAND4BXL U2977 ( .AN(n2241), .B(n2240), .C(n2239), .D(n2238), .Y(n2255) );
  OAI21XL U2978 ( .A0(n2259), .A1(y[74]), .B0(n2258), .Y(n2260) );
  AOI21XL U2979 ( .A0(n2915), .A1(n2261), .B0(n2260), .Y(n2262) );
  AOI21XL U2980 ( .A0(direction[2]), .A1(n2573), .B0(n2586), .Y(n2554) );
  OAI221XL U2981 ( .A0(pri[2]), .A1(n2554), .B0(pri[1]), .B1(n2391), .C0(n2271), .Y(n2272) );
  NOR2X1 U2982 ( .A(n2799), .B(n2838), .Y(n2849) );
  NOR2XL U2983 ( .A(cnt[1]), .B(N2025), .Y(n2275) );
  OAI21XL U2984 ( .A0(n2275), .A1(n2875), .B0(n2790), .Y(n2276) );
  AOI21XL U2985 ( .A0(cs[0]), .A1(n2661), .B0(n2925), .Y(n2278) );
  NAND2XL U2986 ( .A(n2672), .B(n2874), .Y(n1605) );
  NAND2X2 U2987 ( .A(move_out[2]), .B(n2808), .Y(n2292) );
  AOI21XL U2988 ( .A0(n2873), .A1(n2292), .B0(n2810), .Y(n2279) );
  NAND2XL U2989 ( .A(n2672), .B(n2279), .Y(n1602) );
  NAND3X2 U2990 ( .A(n2672), .B(move_out[4]), .C(n2873), .Y(n2293) );
  NOR2X2 U2991 ( .A(n2293), .B(n2296), .Y(n2742) );
  NAND3X2 U2992 ( .A(move_out[3]), .B(n2672), .C(n2926), .Y(n2286) );
  NOR2X2 U2993 ( .A(n2286), .B(n2296), .Y(n2754) );
  AOI22XL U2994 ( .A0(y[26]), .A1(n2754), .B0(y[74]), .B1(n2373), .Y(n2282) );
  NAND2X1 U2995 ( .A(move_out[2]), .B(n2288), .Y(n2290) );
  NOR2X2 U2996 ( .A(n2286), .B(n2290), .Y(n2734) );
  NAND2X1 U2997 ( .A(n2287), .B(move_out[2]), .Y(n2291) );
  NOR2X2 U2998 ( .A(n2286), .B(n2291), .Y(n2737) );
  NAND2X1 U2999 ( .A(move_out[2]), .B(n2807), .Y(n2294) );
  NOR2X2 U3000 ( .A(n2286), .B(n2294), .Y(n2716) );
  NOR2X2 U3001 ( .A(n2286), .B(n2292), .Y(n2746) );
  AOI22XL U3002 ( .A0(y[38]), .A1(n2716), .B0(y[47]), .B1(n2746), .Y(n2280) );
  NOR2X2 U3003 ( .A(n2294), .B(n2295), .Y(n2702) );
  NOR2X2 U3004 ( .A(n2292), .B(n2295), .Y(n2710) );
  NOR2X2 U3005 ( .A(n2290), .B(n2295), .Y(n2706) );
  NOR2X2 U3006 ( .A(n2291), .B(n2295), .Y(n2694) );
  NAND2X1 U3007 ( .A(n2808), .B(n2284), .Y(n2682) );
  INVX1 U3008 ( .A(n2748), .Y(n2632) );
  AOI22XL U3009 ( .A0(y[8]), .A1(n2630), .B0(y[5]), .B1(n2632), .Y(n2285) );
  OAI21XL U3010 ( .A0(n2906), .A1(n2682), .B0(n2285), .Y(n2302) );
  INVX1 U3011 ( .A(n2770), .Y(n2619) );
  INVX1 U3012 ( .A(n2767), .Y(n2576) );
  AOI22XL U3013 ( .A0(n2619), .A1(y[29]), .B0(y[35]), .B1(n2576), .Y(n2300) );
  INVX1 U3014 ( .A(n2763), .Y(n2582) );
  NOR2X2 U3015 ( .A(n2290), .B(n2293), .Y(n2723) );
  AOI22XL U3016 ( .A0(y[32]), .A1(n2582), .B0(y[68]), .B1(n2723), .Y(n2299) );
  NOR2X2 U3017 ( .A(n2291), .B(n2293), .Y(n2726) );
  NOR2X2 U3018 ( .A(n2292), .B(n2293), .Y(n2792) );
  AOI22XL U3019 ( .A0(y[65]), .A1(n2726), .B0(y[71]), .B1(n2792), .Y(n2298) );
  NOR2X2 U3020 ( .A(n2294), .B(n2293), .Y(n2729) );
  NOR2X2 U3021 ( .A(n2296), .B(n2295), .Y(n2698) );
  AOI22XL U3022 ( .A0(y[62]), .A1(n2729), .B0(y[2]), .B1(n2698), .Y(n2297) );
  AOI22XL U3023 ( .A0(x[24]), .A1(n2754), .B0(x[72]), .B1(n2373), .Y(n2311) );
  AOI22XL U3024 ( .A0(x[36]), .A1(n2716), .B0(x[45]), .B1(n2746), .Y(n2309) );
  AOI22XL U3025 ( .A0(x[3]), .A1(n2632), .B0(x[51]), .B1(n2579), .Y(n2312) );
  OAI21XL U3026 ( .A0(n2929), .A1(n2682), .B0(n2312), .Y(n2318) );
  AOI22XL U3027 ( .A0(n2619), .A1(x[27]), .B0(x[33]), .B1(n2576), .Y(n2316) );
  AOI22XL U3028 ( .A0(x[30]), .A1(n2582), .B0(x[66]), .B1(n2723), .Y(n2315) );
  AOI22XL U3029 ( .A0(x[63]), .A1(n2726), .B0(x[69]), .B1(n2792), .Y(n2314) );
  AOI22XL U3030 ( .A0(x[0]), .A1(n2698), .B0(x[60]), .B1(n2729), .Y(n2313) );
  AOI22XL U3031 ( .A0(x[38]), .A1(n2716), .B0(x[47]), .B1(n2746), .Y(n2325) );
  AOI22XL U3032 ( .A0(x[8]), .A1(n2630), .B0(x[5]), .B1(n2632), .Y(n2328) );
  OAI21XL U3033 ( .A0(n2930), .A1(n2682), .B0(n2328), .Y(n2334) );
  AOI22XL U3034 ( .A0(n2619), .A1(x[29]), .B0(x[35]), .B1(n2576), .Y(n2332) );
  AOI22XL U3035 ( .A0(x[32]), .A1(n2582), .B0(x[68]), .B1(n2723), .Y(n2331) );
  AOI22XL U3036 ( .A0(x[65]), .A1(n2726), .B0(x[71]), .B1(n2792), .Y(n2330) );
  AOI22XL U3037 ( .A0(x[62]), .A1(n2729), .B0(x[2]), .B1(n2698), .Y(n2329) );
  AOI22XL U3038 ( .A0(x[25]), .A1(n2754), .B0(x[73]), .B1(n2373), .Y(n2343) );
  AOI22XL U3039 ( .A0(x[37]), .A1(n2716), .B0(x[46]), .B1(n2746), .Y(n2341) );
  AOI22XL U3040 ( .A0(x[7]), .A1(n2630), .B0(x[4]), .B1(n2632), .Y(n2344) );
  OAI21XL U3041 ( .A0(n2931), .A1(n2682), .B0(n2344), .Y(n2350) );
  AOI22XL U3042 ( .A0(n2619), .A1(x[28]), .B0(x[34]), .B1(n2576), .Y(n2348) );
  AOI22XL U3043 ( .A0(x[31]), .A1(n2582), .B0(x[67]), .B1(n2723), .Y(n2347) );
  AOI22XL U3044 ( .A0(x[64]), .A1(n2726), .B0(x[70]), .B1(n2792), .Y(n2346) );
  AOI22XL U3045 ( .A0(x[61]), .A1(n2729), .B0(x[1]), .B1(n2698), .Y(n2345) );
  AOI22XL U3046 ( .A0(y[25]), .A1(n2754), .B0(y[73]), .B1(n2373), .Y(n2359) );
  AOI22XL U3047 ( .A0(y[37]), .A1(n2716), .B0(y[46]), .B1(n2746), .Y(n2357) );
  AOI22XL U3048 ( .A0(y[7]), .A1(n2630), .B0(y[4]), .B1(n2632), .Y(n2360) );
  OAI21XL U3049 ( .A0(n2928), .A1(n2682), .B0(n2360), .Y(n2366) );
  AOI22XL U3050 ( .A0(n2619), .A1(y[28]), .B0(y[34]), .B1(n2576), .Y(n2364) );
  AOI22XL U3051 ( .A0(y[31]), .A1(n2582), .B0(y[67]), .B1(n2723), .Y(n2363) );
  AOI22XL U3052 ( .A0(y[64]), .A1(n2726), .B0(y[70]), .B1(n2792), .Y(n2362) );
  AOI22XL U3053 ( .A0(y[61]), .A1(n2729), .B0(y[1]), .B1(n2698), .Y(n2361) );
  AOI22XL U3054 ( .A0(y[24]), .A1(n2754), .B0(y[72]), .B1(n2373), .Y(n2376) );
  AOI22XL U3055 ( .A0(y[36]), .A1(n2716), .B0(y[45]), .B1(n2746), .Y(n2374) );
  AOI22XL U3056 ( .A0(y[6]), .A1(n2630), .B0(y[3]), .B1(n2632), .Y(n2377) );
  OAI21XL U3057 ( .A0(n2881), .A1(n2682), .B0(n2377), .Y(n2383) );
  AOI22XL U3058 ( .A0(n2619), .A1(y[27]), .B0(y[33]), .B1(n2576), .Y(n2381) );
  AOI22XL U3059 ( .A0(y[30]), .A1(n2582), .B0(y[66]), .B1(n2723), .Y(n2380) );
  AOI22XL U3060 ( .A0(y[63]), .A1(n2726), .B0(y[69]), .B1(n2792), .Y(n2379) );
  AOI22XL U3061 ( .A0(y[60]), .A1(n2729), .B0(y[0]), .B1(n2698), .Y(n2378) );
  INVXL U3062 ( .A(n2391), .Y(n2392) );
  NOR2BX1 U3063 ( .AN(n2401), .B(n2400), .Y(n2507) );
  AOI22XL U3064 ( .A0(n1761), .A1(y[22]), .B0(n1763), .B1(y[16]), .Y(n2398) );
  AOI22XL U3065 ( .A0(n2765), .A1(y[1]), .B0(n1760), .B1(y[4]), .Y(n2397) );
  AOI22XL U3066 ( .A0(n1765), .A1(y[7]), .B0(n1762), .B1(y[13]), .Y(n2396) );
  AOI22XL U3067 ( .A0(n1766), .A1(y[19]), .B0(n1767), .B1(y[10]), .Y(n2395) );
  AOI22XL U3068 ( .A0(n1761), .A1(y[70]), .B0(n1763), .B1(y[64]), .Y(n2405) );
  AOI22XL U3069 ( .A0(n2765), .A1(y[49]), .B0(n1760), .B1(y[52]), .Y(n2404) );
  AOI22XL U3070 ( .A0(n1765), .A1(y[55]), .B0(n1762), .B1(y[61]), .Y(n2403) );
  AOI22XL U3071 ( .A0(n1766), .A1(y[67]), .B0(n1767), .B1(y[58]), .Y(n2402) );
  AOI22XL U3072 ( .A0(n1761), .A1(y[46]), .B0(n1763), .B1(y[40]), .Y(n2411) );
  AOI22XL U3073 ( .A0(n2765), .A1(y[25]), .B0(n1760), .B1(y[28]), .Y(n2410) );
  AOI22XL U3074 ( .A0(y[31]), .A1(n1765), .B0(y[37]), .B1(n1762), .Y(n2409) );
  AOI22XL U3075 ( .A0(n1766), .A1(y[43]), .B0(y[34]), .B1(n1767), .Y(n2408) );
  OAI21XL U3076 ( .A0(n2910), .A1(n2488), .B0(n2414), .Y(n2415) );
  AOI22XL U3077 ( .A0(n1761), .A1(y[21]), .B0(n1763), .B1(y[15]), .Y(n2420) );
  AOI22XL U3078 ( .A0(n2765), .A1(y[0]), .B0(n1760), .B1(y[3]), .Y(n2419) );
  AOI22XL U3079 ( .A0(n1765), .A1(y[6]), .B0(n1762), .B1(y[12]), .Y(n2418) );
  AOI22XL U3080 ( .A0(n1766), .A1(y[18]), .B0(n1767), .B1(y[9]), .Y(n2417) );
  AOI22XL U3081 ( .A0(n1761), .A1(y[45]), .B0(n1763), .B1(y[39]), .Y(n2425) );
  AOI22XL U3082 ( .A0(n2765), .A1(y[24]), .B0(n1760), .B1(y[27]), .Y(n2424) );
  AOI22XL U3083 ( .A0(n1765), .A1(y[30]), .B0(n1762), .B1(y[36]), .Y(n2423) );
  AOI22XL U3084 ( .A0(n1766), .A1(y[42]), .B0(n1767), .B1(y[33]), .Y(n2422) );
  AOI22XL U3085 ( .A0(n1761), .A1(y[69]), .B0(n1763), .B1(y[63]), .Y(n2429) );
  AOI22XL U3086 ( .A0(n2765), .A1(y[48]), .B0(n1760), .B1(y[51]), .Y(n2428) );
  AOI22XL U3087 ( .A0(n1765), .A1(y[54]), .B0(n1762), .B1(y[60]), .Y(n2427) );
  AOI22XL U3088 ( .A0(n1766), .A1(y[66]), .B0(n1767), .B1(y[57]), .Y(n2426) );
  AOI22XL U3089 ( .A0(n1761), .A1(y[23]), .B0(n1763), .B1(y[17]), .Y(n2437) );
  AOI22XL U3090 ( .A0(n2765), .A1(y[2]), .B0(n1760), .B1(y[5]), .Y(n2436) );
  AOI22XL U3091 ( .A0(n1765), .A1(y[8]), .B0(n1762), .B1(y[14]), .Y(n2435) );
  AOI22XL U3092 ( .A0(n1766), .A1(y[20]), .B0(n1767), .B1(y[11]), .Y(n2434) );
  AOI22XL U3093 ( .A0(n1761), .A1(y[71]), .B0(n1763), .B1(y[65]), .Y(n2441) );
  AOI22XL U3094 ( .A0(n2765), .A1(y[50]), .B0(n1760), .B1(y[53]), .Y(n2440) );
  AOI22XL U3095 ( .A0(n1765), .A1(y[56]), .B0(n1762), .B1(y[62]), .Y(n2439) );
  AOI22XL U3096 ( .A0(n1766), .A1(y[68]), .B0(n1767), .B1(y[59]), .Y(n2438) );
  AOI22XL U3097 ( .A0(n1761), .A1(y[47]), .B0(n1763), .B1(y[41]), .Y(n2445) );
  AOI22XL U3098 ( .A0(n2765), .A1(y[26]), .B0(n1760), .B1(y[29]), .Y(n2444) );
  AOI22XL U3099 ( .A0(n1765), .A1(y[32]), .B0(n1762), .B1(y[38]), .Y(n2443) );
  AOI22XL U3100 ( .A0(n1766), .A1(y[44]), .B0(n1767), .B1(y[35]), .Y(n2442) );
  OAI21XL U3101 ( .A0(n2908), .A1(n2488), .B0(n2448), .Y(n2449) );
  INVXL U3102 ( .A(n2527), .Y(n2454) );
  OAI21XL U3103 ( .A0(n2530), .A1(n2454), .B0(n2453), .Y(n2455) );
  AOI22XL U3104 ( .A0(n1761), .A1(x[71]), .B0(n1763), .B1(x[65]), .Y(n2459) );
  AOI22XL U3105 ( .A0(n2765), .A1(x[50]), .B0(n1760), .B1(x[53]), .Y(n2458) );
  AOI22XL U3106 ( .A0(n1765), .A1(x[56]), .B0(n1762), .B1(x[62]), .Y(n2457) );
  AOI22XL U3107 ( .A0(n1766), .A1(x[68]), .B0(n1767), .B1(x[59]), .Y(n2456) );
  AOI22XL U3108 ( .A0(n1761), .A1(x[47]), .B0(n1763), .B1(x[41]), .Y(n2464) );
  AOI22XL U3109 ( .A0(n2785), .A1(x[26]), .B0(n1760), .B1(x[29]), .Y(n2463) );
  AOI22XL U3110 ( .A0(n1765), .A1(x[32]), .B0(n1762), .B1(x[38]), .Y(n2462) );
  AOI22XL U3111 ( .A0(n1766), .A1(x[44]), .B0(n1767), .B1(x[35]), .Y(n2461) );
  AOI22XL U3112 ( .A0(n1761), .A1(x[23]), .B0(n1763), .B1(x[17]), .Y(n2468) );
  AOI22XL U3113 ( .A0(n2785), .A1(x[2]), .B0(n1760), .B1(x[5]), .Y(n2467) );
  AOI22XL U3114 ( .A0(n1765), .A1(x[8]), .B0(n1762), .B1(x[14]), .Y(n2466) );
  AOI22XL U3115 ( .A0(n1766), .A1(x[20]), .B0(n1767), .B1(x[11]), .Y(n2465) );
  AOI22XL U3116 ( .A0(n1761), .A1(x[45]), .B0(n1763), .B1(x[39]), .Y(n2476) );
  AOI22XL U3117 ( .A0(n2785), .A1(x[24]), .B0(n1760), .B1(x[27]), .Y(n2475) );
  AOI22XL U3118 ( .A0(n1765), .A1(x[30]), .B0(n1762), .B1(x[36]), .Y(n2474) );
  AOI22XL U3119 ( .A0(n1766), .A1(x[42]), .B0(n1767), .B1(x[33]), .Y(n2473) );
  AOI22XL U3120 ( .A0(n1761), .A1(x[69]), .B0(n1763), .B1(x[63]), .Y(n2480) );
  AOI22XL U3121 ( .A0(n1859), .A1(x[48]), .B0(n1760), .B1(x[51]), .Y(n2479) );
  AOI22XL U3122 ( .A0(n1765), .A1(x[54]), .B0(n1762), .B1(x[60]), .Y(n2478) );
  AOI22XL U3123 ( .A0(n1766), .A1(x[66]), .B0(n1767), .B1(x[57]), .Y(n2477) );
  AOI22XL U3124 ( .A0(n1761), .A1(x[21]), .B0(n1763), .B1(x[15]), .Y(n2484) );
  AOI22XL U3125 ( .A0(n1859), .A1(x[0]), .B0(n1760), .B1(x[3]), .Y(n2483) );
  AOI22XL U3126 ( .A0(n1765), .A1(x[6]), .B0(n1762), .B1(x[12]), .Y(n2482) );
  AOI22XL U3127 ( .A0(n1766), .A1(x[18]), .B0(n1767), .B1(x[9]), .Y(n2481) );
  OAI21XL U3128 ( .A0(n2911), .A1(n2488), .B0(n2487), .Y(n2489) );
  AOI22XL U3129 ( .A0(n1761), .A1(x[70]), .B0(n1763), .B1(x[64]), .Y(n2494) );
  AOI22XL U3130 ( .A0(n2785), .A1(x[49]), .B0(n1760), .B1(x[52]), .Y(n2493) );
  AOI22XL U3131 ( .A0(n1765), .A1(x[55]), .B0(n1762), .B1(x[61]), .Y(n2492) );
  AOI22XL U3132 ( .A0(n1766), .A1(x[67]), .B0(n1767), .B1(x[58]), .Y(n2491) );
  AOI22XL U3133 ( .A0(n1761), .A1(x[46]), .B0(n1763), .B1(x[40]), .Y(n2501) );
  AOI22XL U3134 ( .A0(n2785), .A1(x[25]), .B0(n1760), .B1(x[28]), .Y(n2500) );
  AOI22XL U3135 ( .A0(n1765), .A1(x[31]), .B0(n1762), .B1(x[37]), .Y(n2499) );
  AOI22XL U3136 ( .A0(n1766), .A1(x[43]), .B0(n1767), .B1(x[34]), .Y(n2498) );
  AOI22XL U3137 ( .A0(n1761), .A1(x[22]), .B0(n1763), .B1(x[16]), .Y(n2505) );
  AOI22XL U3138 ( .A0(n2785), .A1(x[1]), .B0(n1760), .B1(x[4]), .Y(n2504) );
  AOI22XL U3139 ( .A0(n1765), .A1(x[7]), .B0(n1762), .B1(x[13]), .Y(n2503) );
  AOI22XL U3140 ( .A0(n1766), .A1(x[19]), .B0(n1767), .B1(x[10]), .Y(n2502) );
  AOI21XL U3141 ( .A0(n2513), .A1(n2512), .B0(n2520), .Y(n2541) );
  OAI21XL U3142 ( .A0(n2515), .A1(n2514), .B0(n2516), .Y(n2539) );
  CMPR32X1 U3143 ( .A(n2518), .B(n2517), .C(n2516), .CO(n2452), .S(n2543) );
  CMPR32X1 U3144 ( .A(n2521), .B(n2520), .C(n2519), .CO(n2522), .S(n2542) );
  CMPR32X1 U3145 ( .A(n2524), .B(n2523), .C(n2522), .CO(n2537), .S(n2538) );
  OAI21XL U3146 ( .A0(n2530), .A1(n2529), .B0(n2527), .Y(n2528) );
  NAND4BXL U3147 ( .AN(n2542), .B(n2541), .C(n2540), .D(n2539), .Y(n2546) );
  OAI211X1 U3148 ( .A0(n2545), .A1(n2556), .B0(n2557), .C0(n2544), .Y(n2850)
         );
  AOI21XL U3149 ( .A0(n2850), .A1(n2563), .B0(n2638), .Y(n2548) );
  OAI21XL U3150 ( .A0(n2850), .A1(n2563), .B0(n2548), .Y(n2550) );
  OAI21XL U3151 ( .A0(n2559), .A1(n2558), .B0(n2557), .Y(n2560) );
  AOI21XL U3152 ( .A0(n2566), .A1(n2565), .B0(n2638), .Y(n2564) );
  OAI21XL U3153 ( .A0(n2566), .A1(n2565), .B0(n2564), .Y(n2567) );
  NOR2X4 U3154 ( .A(n2713), .B(n2628), .Y(n2620) );
  AOI21X2 U3155 ( .A0(n1763), .A1(n2620), .B0(n2746), .Y(n2612) );
  NOR2X2 U3156 ( .A(n2732), .B(n2621), .Y(n2611) );
  NOR2X4 U3157 ( .A(n2718), .B(n2628), .Y(n2580) );
  AOI21X2 U3158 ( .A0(n1762), .A1(n2580), .B0(n2723), .Y(n2618) );
  NOR2X2 U3159 ( .A(n2735), .B(n2581), .Y(n2617) );
  AOI21X2 U3160 ( .A0(n1760), .A1(n2580), .B0(n2574), .Y(n2602) );
  NOR2X2 U3161 ( .A(n2578), .B(n2581), .Y(n2601) );
  AOI21X2 U3162 ( .A0(n1762), .A1(n2620), .B0(n2734), .Y(n2604) );
  NOR2X2 U3163 ( .A(n2735), .B(n2621), .Y(n2603) );
  AOI21X2 U3164 ( .A0(n1763), .A1(n2580), .B0(n2792), .Y(n2616) );
  NOR2X2 U3165 ( .A(n2732), .B(n2581), .Y(n2615) );
  AOI21X2 U3166 ( .A0(n2765), .A1(n2580), .B0(n2575), .Y(n2610) );
  NOR2X2 U3167 ( .A(n2780), .B(n2581), .Y(n2609) );
  AOI21X2 U3168 ( .A0(n2738), .A1(n2580), .B0(n2726), .Y(n2614) );
  NOR2X2 U3169 ( .A(n2727), .B(n2581), .Y(n2613) );
  AOI21X2 U3170 ( .A0(n1760), .A1(n2620), .B0(n2576), .Y(n2596) );
  NOR2X2 U3171 ( .A(n2578), .B(n2621), .Y(n2595) );
  AOI21X2 U3172 ( .A0(n2738), .A1(n2620), .B0(n2737), .Y(n2600) );
  NOR2X2 U3173 ( .A(n2727), .B(n2621), .Y(n2599) );
  AOI21X2 U3174 ( .A0(n1761), .A1(n2580), .B0(n2579), .Y(n2606) );
  NOR2X2 U3175 ( .A(n2752), .B(n2581), .Y(n2605) );
  AOI21X2 U3176 ( .A0(n1765), .A1(n2580), .B0(n2729), .Y(n2608) );
  NOR2X2 U3177 ( .A(n2776), .B(n2581), .Y(n2607) );
  AOI21X2 U3178 ( .A0(n2765), .A1(n2620), .B0(n2582), .Y(n2598) );
  NOR2X2 U3179 ( .A(n2780), .B(n2621), .Y(n2597) );
  AOI21X2 U3180 ( .A0(n1765), .A1(n2620), .B0(n2716), .Y(n2594) );
  NOR2X2 U3181 ( .A(n2776), .B(n2621), .Y(n2593) );
  AND2X2 U3182 ( .A(n2588), .B(n2591), .Y(n2664) );
  AND2X2 U3183 ( .A(n2589), .B(n2591), .Y(n2665) );
  AND2X2 U3184 ( .A(n2590), .B(n2591), .Y(n2668) );
  AND2X2 U3185 ( .A(n2592), .B(n2591), .Y(n2666) );
  AOI21X2 U3186 ( .A0(n1761), .A1(n2620), .B0(n2619), .Y(n2627) );
  NOR2X2 U3187 ( .A(n2752), .B(n2621), .Y(n2626) );
  AOI21X2 U3188 ( .A0(n2662), .A1(n2707), .B0(n2706), .Y(n2656) );
  NOR2X2 U3189 ( .A(n1769), .B(n2629), .Y(n2655) );
  AOI21X2 U3190 ( .A0(n2662), .A1(n2743), .B0(n2742), .Y(n2648) );
  AOI21X2 U3191 ( .A0(n2662), .A1(n2761), .B0(n2630), .Y(n2652) );
  NOR2X2 U3192 ( .A(n1769), .B(n2631), .Y(n2651) );
  AOI21X2 U3193 ( .A0(n2662), .A1(n2750), .B0(n2632), .Y(n2644) );
  NOR2X2 U3194 ( .A(n1769), .B(n2633), .Y(n2643) );
  AOI21X2 U3195 ( .A0(n2662), .A1(n2703), .B0(n2702), .Y(n2650) );
  NOR2X2 U3196 ( .A(n1769), .B(n2634), .Y(n2649) );
  AOI21X2 U3197 ( .A0(n2662), .A1(n2699), .B0(n2698), .Y(n2642) );
  NOR2X2 U3198 ( .A(n1769), .B(n2635), .Y(n2641) );
  AOI21X2 U3199 ( .A0(n2662), .A1(n2695), .B0(n2694), .Y(n2646) );
  NOR2X2 U3200 ( .A(n1769), .B(n2636), .Y(n2645) );
  AOI21X2 U3201 ( .A0(n2662), .A1(n2711), .B0(n2710), .Y(n2654) );
  NOR2X2 U3202 ( .A(n1769), .B(n2637), .Y(n2653) );
  AOI21X2 U3203 ( .A0(n2662), .A1(n2755), .B0(n2754), .Y(n2658) );
  AOI21X2 U3204 ( .A0(n2662), .A1(n2684), .B0(n2639), .Y(n2660) );
  NOR2X2 U3205 ( .A(n1769), .B(n2640), .Y(n2659) );
  AOI31X4 U3206 ( .A0(n2674), .A1(n1766), .A2(n2662), .B0(n2673), .Y(n2669) );
  NOR2X2 U3207 ( .A(n1769), .B(n2663), .Y(n2667) );
  NOR2X2 U3208 ( .A(n2672), .B(n2671), .Y(n2801) );
  OAI21XL U3209 ( .A0(n1849), .A1(n2797), .B0(n1595), .Y(n2676) );
  AOI21XL U3210 ( .A0(n2801), .A1(in_x[1]), .B0(n2676), .Y(n2677) );
  OAI21XL U3211 ( .A0(n2758), .A1(n2776), .B0(n2682), .Y(n2683) );
  NOR2X2 U3212 ( .A(n2719), .B(n2713), .Y(n2773) );
  NOR2X2 U3213 ( .A(n2719), .B(n2718), .Y(n2793) );
  OAI21XL U3214 ( .A0(n2758), .A1(n2780), .B0(n2748), .Y(n2749) );
  OAI21XL U3215 ( .A0(n2758), .A1(n2578), .B0(n2757), .Y(n2759) );
  OAI21XL U3216 ( .A0(n2771), .A1(n2578), .B0(n2763), .Y(n2764) );
  OAI21XL U3217 ( .A0(n2771), .A1(n2776), .B0(n2767), .Y(n2768) );
  OAI21XL U3218 ( .A0(n2780), .A1(n2771), .B0(n2770), .Y(n2772) );
  OAI21XL U3219 ( .A0(n2789), .A1(n2776), .B0(n2775), .Y(n2777) );
  OAI21XL U3220 ( .A0(n2780), .A1(n2789), .B0(n2779), .Y(n2781) );
  OAI21XL U3221 ( .A0(n2789), .A1(n2578), .B0(n2783), .Y(n2784) );
  AOI21XL U3222 ( .A0(move_out[4]), .A1(n2810), .B0(n1595), .Y(n2809) );
  OAI21XL U3223 ( .A0(move_out[4]), .A1(n2810), .B0(n2809), .Y(n1601) );
  INVXL U3224 ( .A(n2840), .Y(n2839) );
  OAI21XL U3225 ( .A0(n2842), .A1(n2846), .B0(n2841), .Y(n2843) );
  AOI21XL U3226 ( .A0(cnt[4]), .A1(n2849), .B0(n2843), .Y(n1593) );
  OAI21XL U3227 ( .A0(cnt[1]), .A1(N2025), .B0(n2844), .Y(n2845) );
  AOI21XL U3228 ( .A0(cnt[1]), .A1(n2849), .B0(n2848), .Y(n1591) );
  OAI21XL U3229 ( .A0(n2858), .A1(n2857), .B0(n2856), .Y(n2859) );
  AOI21XL U3230 ( .A0(direction[0]), .A1(n2860), .B0(n2859), .Y(n1585) );
endmodule


